
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-32.95,39.6893,61.95,-63.2229</PageViewport>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>14.5,-13</position>
<gparam>LABEL_TEXT Go to https://cedar.to/vjyQw7 to download the latest version!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_LABEL</type>
<position>14.5,-9.5</position>
<gparam>LABEL_TEXT Error: This file was made with a newer version of Cedar Logic!</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate></page 0>
</circuit>
<throw_away></throw_away>

	<version>2.3.6 | 2021-11-12 10:52:37</version><circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-164.331,64.2856,274.593,-147.945</PageViewport>
<gate>
<ID>73</ID>
<type>BE_JKFF_LOW_NT</type>
<position>18,-110</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>52 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>9</ID>
<type>DA_FROM</type>
<position>34,-24</position>
<input>
<ID>IN_0</ID>8 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>65</ID>
<type>DA_FROM</type>
<position>2,-86</position>
<input>
<ID>IN_0</ID>43 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>1</ID>
<type>BE_JKFF_LOW_NT</type>
<position>50,-17</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>3 </output>
<input>
<ID>clock</ID>1 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>74</ID>
<type>BE_JKFF_LOW_NT</type>
<position>7.5,-110</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>53 </output>
<input>
<ID>clock</ID>52 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>10</ID>
<type>DA_FROM</type>
<position>24,-24</position>
<input>
<ID>IN_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>2</ID>
<type>BE_JKFF_LOW_NT</type>
<position>39.5,-17</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>8 </output>
<input>
<ID>clock</ID>3 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>3</ID>
<type>BB_CLOCK</type>
<position>54.5,-23.5</position>
<output>
<ID>CLK</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>4</ID>
<type>BE_JKFF_LOW_NT</type>
<position>29,-17</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>4 </output>
<input>
<ID>clock</ID>8 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>5</ID>
<type>BE_JKFF_LOW_NT</type>
<position>18.5,-17</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>5 </output>
<input>
<ID>clock</ID>4 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>70</ID>
<type>BE_JKFF_LOW_NT</type>
<position>49.5,-110</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>50 </output>
<input>
<ID>clock</ID>48 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>6</ID>
<type>BE_JKFF_LOW_NT</type>
<position>8,-17</position>
<input>
<ID>J</ID>2 </input>
<input>
<ID>K</ID>2 </input>
<output>
<ID>Q</ID>6 </output>
<input>
<ID>clock</ID>5 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>11</ID>
<type>DA_FROM</type>
<position>13,-24</position>
<input>
<ID>IN_0</ID>5 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>12</ID>
<type>DA_FROM</type>
<position>3,-24</position>
<input>
<ID>IN_0</ID>6 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>77</ID>
<type>BB_CLOCK</type>
<position>54.5,-116.5</position>
<output>
<ID>CLK</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>13</ID>
<type>GA_LED</type>
<position>175.5,-80</position>
<input>
<ID>N_in0</ID>23 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BE_JKFF_LOW_NT</type>
<position>49.5,-50</position>
<input>
<ID>J</ID>29 </input>
<input>
<ID>K</ID>29 </input>
<output>
<ID>Q</ID>30 </output>
<input>
<ID>clock</ID>28 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>21</ID>
<type>BE_JKFF_LOW_NT</type>
<position>39,-50</position>
<input>
<ID>J</ID>29 </input>
<input>
<ID>K</ID>29 </input>
<output>
<ID>Q</ID>35 </output>
<input>
<ID>clock</ID>30 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>23</ID>
<type>BE_JKFF_LOW_NT</type>
<position>28.5,-50</position>
<input>
<ID>J</ID>29 </input>
<input>
<ID>K</ID>29 </input>
<output>
<ID>Q</ID>31 </output>
<input>
<ID>clock</ID>35 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>25</ID>
<type>BE_JKFF_LOW_NT</type>
<position>7.5,-50</position>
<input>
<ID>J</ID>29 </input>
<input>
<ID>K</ID>29 </input>
<output>
<ID>Q</ID>33 </output>
<input>
<ID>clock</ID>32 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>29</ID>
<type>BB_CLOCK</type>
<position>53,-56.5</position>
<output>
<ID>CLK</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>31</ID>
<type>DA_FROM</type>
<position>23.5,-57</position>
<input>
<ID>IN_0</ID>31 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>33</ID>
<type>DA_FROM</type>
<position>12.5,-57</position>
<input>
<ID>IN_0</ID>32 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>34</ID>
<type>AE_DFF_LOW</type>
<position>142,-63.5</position>
<input>
<ID>IN_0</ID>164 </input>
<output>
<ID>OUT_0</ID>19 </output>
<input>
<ID>clear</ID>21 </input>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>35</ID>
<type>DA_FROM</type>
<position>2.5,-57</position>
<input>
<ID>IN_0</ID>33 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>36</ID>
<type>AE_DFF_LOW</type>
<position>142.5,-23.5</position>
<input>
<ID>IN_0</ID>156 </input>
<output>
<ID>OUT_0</ID>22 </output>
<input>
<ID>clear</ID>21 </input>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>166</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-26.5,-17</position>
<input>
<ID>J</ID>127 </input>
<input>
<ID>K</ID>127 </input>
<output>
<ID>Q</ID>132 </output>
<input>
<ID>clock</ID>128 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>38</ID>
<type>AE_DFF_LOW</type>
<position>142.5,-47</position>
<input>
<ID>IN_0</ID>163 </input>
<output>
<ID>OUT_0</ID>20 </output>
<input>
<ID>clear</ID>21 </input>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>168</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-37,-17</position>
<input>
<ID>J</ID>127 </input>
<input>
<ID>K</ID>127 </input>
<output>
<ID>Q</ID>129 </output>
<input>
<ID>clock</ID>132 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>174.5,-61</position>
<input>
<ID>N_in0</ID>19 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-47.5,-17</position>
<input>
<ID>J</ID>127 </input>
<input>
<ID>K</ID>127 </input>
<output>
<ID>Q</ID>130 </output>
<input>
<ID>clock</ID>129 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>41</ID>
<type>GA_LED</type>
<position>173,-17.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-58,-17</position>
<input>
<ID>J</ID>127 </input>
<input>
<ID>K</ID>127 </input>
<output>
<ID>Q</ID>131 </output>
<input>
<ID>clock</ID>130 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>42</ID>
<type>BE_JKFF_LOW_NT</type>
<position>49,-79</position>
<input>
<ID>J</ID>39 </input>
<input>
<ID>K</ID>39 </input>
<output>
<ID>Q</ID>40 </output>
<input>
<ID>clock</ID>38 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>171</ID>
<type>DA_FROM</type>
<position>-32,-24</position>
<input>
<ID>IN_0</ID>132 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>43</ID>
<type>GA_LED</type>
<position>172,-37.5</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>DA_FROM</type>
<position>-53,-24</position>
<input>
<ID>IN_0</ID>130 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>45</ID>
<type>AE_DFF_LOW</type>
<position>141.5,-82</position>
<input>
<ID>IN_0</ID>165 </input>
<output>
<ID>OUT_0</ID>23 </output>
<input>
<ID>clear</ID>21 </input>
<input>
<ID>clock</ID>18 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>52</ID>
<type>BE_JKFF_LOW_NT</type>
<position>18,-50</position>
<input>
<ID>J</ID>29 </input>
<input>
<ID>K</ID>29 </input>
<output>
<ID>Q</ID>32 </output>
<input>
<ID>clock</ID>31 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>54</ID>
<type>DA_FROM</type>
<position>33.5,-57</position>
<input>
<ID>IN_0</ID>35 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>56</ID>
<type>BE_JKFF_LOW_NT</type>
<position>38.5,-79</position>
<input>
<ID>J</ID>39 </input>
<input>
<ID>K</ID>39 </input>
<output>
<ID>Q</ID>45 </output>
<input>
<ID>clock</ID>40 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>57</ID>
<type>BE_JKFF_LOW_NT</type>
<position>28,-79</position>
<input>
<ID>J</ID>39 </input>
<input>
<ID>K</ID>39 </input>
<output>
<ID>Q</ID>41 </output>
<input>
<ID>clock</ID>45 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>58</ID>
<type>BE_JKFF_LOW_NT</type>
<position>17.5,-79</position>
<input>
<ID>J</ID>39 </input>
<input>
<ID>K</ID>39 </input>
<output>
<ID>Q</ID>42 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>BE_JKFF_LOW_NT</type>
<position>7,-79</position>
<input>
<ID>J</ID>39 </input>
<input>
<ID>K</ID>39 </input>
<output>
<ID>Q</ID>43 </output>
<input>
<ID>clock</ID>42 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>61</ID>
<type>BB_CLOCK</type>
<position>54,-85.5</position>
<output>
<ID>CLK</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>62</ID>
<type>DA_FROM</type>
<position>33,-86</position>
<input>
<ID>IN_0</ID>45 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>63</ID>
<type>DA_FROM</type>
<position>23,-86</position>
<input>
<ID>IN_0</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>64</ID>
<type>DA_FROM</type>
<position>12,-86</position>
<input>
<ID>IN_0</ID>42 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>71</ID>
<type>BE_JKFF_LOW_NT</type>
<position>39,-110</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>55 </output>
<input>
<ID>clock</ID>50 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>72</ID>
<type>BE_JKFF_LOW_NT</type>
<position>28.5,-110</position>
<input>
<ID>J</ID>49 </input>
<input>
<ID>K</ID>49 </input>
<output>
<ID>Q</ID>51 </output>
<input>
<ID>clock</ID>55 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>78</ID>
<type>DA_FROM</type>
<position>33.5,-117</position>
<input>
<ID>IN_0</ID>55 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>79</ID>
<type>DA_FROM</type>
<position>23.5,-117</position>
<input>
<ID>IN_0</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>80</ID>
<type>DA_FROM</type>
<position>12.5,-117</position>
<input>
<ID>IN_0</ID>52 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>81</ID>
<type>DA_FROM</type>
<position>2.5,-117</position>
<input>
<ID>IN_0</ID>53 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>160</ID>
<type>BB_CLOCK</type>
<position>128,-30.5</position>
<output>
<ID>CLK</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>165</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-16,-17</position>
<input>
<ID>J</ID>127 </input>
<input>
<ID>K</ID>127 </input>
<output>
<ID>Q</ID>128 </output>
<input>
<ID>clock</ID>126 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>167</ID>
<type>BB_CLOCK</type>
<position>-11.5,-23.5</position>
<output>
<ID>CLK</ID>126 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>172</ID>
<type>DA_FROM</type>
<position>-42,-24</position>
<input>
<ID>IN_0</ID>129 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>174</ID>
<type>DA_FROM</type>
<position>-63,-24</position>
<input>
<ID>IN_0</ID>131 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>175</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-16.5,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>135 </output>
<input>
<ID>clock</ID>133 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>176</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-27,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>139 </output>
<input>
<ID>clock</ID>135 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>177</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-37.5,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>136 </output>
<input>
<ID>clock</ID>139 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>178</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-58.5,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>138 </output>
<input>
<ID>clock</ID>137 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>179</ID>
<type>BB_CLOCK</type>
<position>-13,-56.5</position>
<output>
<ID>CLK</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>180</ID>
<type>DA_FROM</type>
<position>-42.5,-57</position>
<input>
<ID>IN_0</ID>136 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F1</lparam></gate>
<gate>
<ID>181</ID>
<type>DA_FROM</type>
<position>-53.5,-57</position>
<input>
<ID>IN_0</ID>137 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G1</lparam></gate>
<gate>
<ID>182</ID>
<type>DA_FROM</type>
<position>-63.5,-57</position>
<input>
<ID>IN_0</ID>138 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H1</lparam></gate>
<gate>
<ID>183</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-17,-79</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>141 </input>
<output>
<ID>Q</ID>142 </output>
<input>
<ID>clock</ID>140 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>184</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-48,-50</position>
<input>
<ID>J</ID>134 </input>
<input>
<ID>K</ID>134 </input>
<output>
<ID>Q</ID>137 </output>
<input>
<ID>clock</ID>136 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>185</ID>
<type>DA_FROM</type>
<position>-32.5,-57</position>
<input>
<ID>IN_0</ID>139 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E1</lparam></gate>
<gate>
<ID>186</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-27.5,-79</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>141 </input>
<output>
<ID>Q</ID>146 </output>
<input>
<ID>clock</ID>142 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>187</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-38,-79</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>141 </input>
<output>
<ID>Q</ID>143 </output>
<input>
<ID>clock</ID>146 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>188</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-48.5,-79</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>141 </input>
<output>
<ID>Q</ID>144 </output>
<input>
<ID>clock</ID>143 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>189</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-59,-79</position>
<input>
<ID>J</ID>141 </input>
<input>
<ID>K</ID>141 </input>
<output>
<ID>Q</ID>145 </output>
<input>
<ID>clock</ID>144 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>190</ID>
<type>BB_CLOCK</type>
<position>-12,-85.5</position>
<output>
<ID>CLK</ID>140 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>191</ID>
<type>DA_FROM</type>
<position>-33,-86</position>
<input>
<ID>IN_0</ID>146 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E2</lparam></gate>
<gate>
<ID>192</ID>
<type>DA_FROM</type>
<position>-43,-86</position>
<input>
<ID>IN_0</ID>143 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F2</lparam></gate>
<gate>
<ID>193</ID>
<type>DA_FROM</type>
<position>-54,-86</position>
<input>
<ID>IN_0</ID>144 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G2</lparam></gate>
<gate>
<ID>194</ID>
<type>DA_FROM</type>
<position>-64,-86</position>
<input>
<ID>IN_0</ID>145 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H2</lparam></gate>
<gate>
<ID>195</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-16.5,-110</position>
<input>
<ID>J</ID>148 </input>
<input>
<ID>K</ID>148 </input>
<output>
<ID>Q</ID>149 </output>
<input>
<ID>clock</ID>147 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>196</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-27,-110</position>
<input>
<ID>J</ID>148 </input>
<input>
<ID>K</ID>148 </input>
<output>
<ID>Q</ID>153 </output>
<input>
<ID>clock</ID>149 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>197</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-37.5,-110</position>
<input>
<ID>J</ID>148 </input>
<input>
<ID>K</ID>148 </input>
<output>
<ID>Q</ID>150 </output>
<input>
<ID>clock</ID>153 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>198</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-48,-110</position>
<input>
<ID>J</ID>148 </input>
<input>
<ID>K</ID>148 </input>
<output>
<ID>Q</ID>151 </output>
<input>
<ID>clock</ID>150 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>199</ID>
<type>BE_JKFF_LOW_NT</type>
<position>-58.5,-110</position>
<input>
<ID>J</ID>148 </input>
<input>
<ID>K</ID>148 </input>
<output>
<ID>Q</ID>152 </output>
<input>
<ID>clock</ID>151 </input>
<gparam>angle 180</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>200</ID>
<type>BB_CLOCK</type>
<position>-11.5,-116.5</position>
<output>
<ID>CLK</ID>147 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 5</lparam></gate>
<gate>
<ID>201</ID>
<type>DA_FROM</type>
<position>-32.5,-117</position>
<input>
<ID>IN_0</ID>153 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID E3</lparam></gate>
<gate>
<ID>202</ID>
<type>DA_FROM</type>
<position>-42.5,-117</position>
<input>
<ID>IN_0</ID>150 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID F3</lparam></gate>
<gate>
<ID>203</ID>
<type>DA_FROM</type>
<position>-53.5,-117</position>
<input>
<ID>IN_0</ID>151 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID G3</lparam></gate>
<gate>
<ID>204</ID>
<type>DA_FROM</type>
<position>-63.5,-117</position>
<input>
<ID>IN_0</ID>152 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID H3</lparam></gate>
<gate>
<ID>212</ID>
<type>AA_AND4</type>
<position>79,-16.5</position>
<input>
<ID>IN_0</ID>172 </input>
<input>
<ID>IN_1</ID>173 </input>
<input>
<ID>IN_2</ID>174 </input>
<input>
<ID>IN_3</ID>175 </input>
<output>
<ID>OUT</ID>154 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>214</ID>
<type>AA_AND3</type>
<position>91.5,-21</position>
<input>
<ID>IN_0</ID>154 </input>
<input>
<ID>IN_1</ID>182 </input>
<input>
<ID>IN_2</ID>155 </input>
<output>
<ID>OUT</ID>156 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>216</ID>
<type>AA_AND4</type>
<position>78.5,-29</position>
<input>
<ID>IN_0</ID>179 </input>
<input>
<ID>IN_1</ID>177 </input>
<input>
<ID>IN_2</ID>178 </input>
<input>
<ID>IN_3</ID>181 </input>
<output>
<ID>OUT</ID>155 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>217</ID>
<type>AA_AND4</type>
<position>79,-40.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>57 </input>
<input>
<ID>IN_2</ID>59 </input>
<input>
<ID>IN_3</ID>60 </input>
<output>
<ID>OUT</ID>157 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>218</ID>
<type>AA_AND3</type>
<position>91.5,-45</position>
<input>
<ID>IN_0</ID>157 </input>
<input>
<ID>IN_1</ID>27 </input>
<input>
<ID>IN_2</ID>158 </input>
<output>
<ID>OUT</ID>163 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND4</type>
<position>78.5,-53</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>62 </input>
<input>
<ID>IN_2</ID>63 </input>
<input>
<ID>IN_3</ID>64 </input>
<output>
<ID>OUT</ID>158 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND4</type>
<position>79,-65</position>
<input>
<ID>IN_0</ID>99 </input>
<input>
<ID>IN_1</ID>98 </input>
<input>
<ID>IN_2</ID>97 </input>
<input>
<ID>IN_3</ID>96 </input>
<output>
<ID>OUT</ID>159 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND3</type>
<position>91.5,-69.5</position>
<input>
<ID>IN_0</ID>159 </input>
<input>
<ID>IN_1</ID>81 </input>
<input>
<ID>IN_2</ID>160 </input>
<output>
<ID>OUT</ID>164 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_AND4</type>
<position>78.5,-77.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>94 </input>
<input>
<ID>IN_2</ID>93 </input>
<input>
<ID>IN_3</ID>92 </input>
<output>
<ID>OUT</ID>160 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_AND4</type>
<position>78.5,-89.5</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>108 </input>
<input>
<ID>IN_2</ID>176 </input>
<input>
<ID>IN_3</ID>190 </input>
<output>
<ID>OUT</ID>161 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>224</ID>
<type>AA_AND3</type>
<position>91,-94</position>
<input>
<ID>IN_0</ID>161 </input>
<input>
<ID>IN_1</ID>82 </input>
<input>
<ID>IN_2</ID>162 </input>
<output>
<ID>OUT</ID>165 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>225</ID>
<type>AA_AND4</type>
<position>78,-102</position>
<input>
<ID>IN_0</ID>103 </input>
<input>
<ID>IN_1</ID>110 </input>
<input>
<ID>IN_2</ID>193 </input>
<input>
<ID>IN_3</ID>192 </input>
<output>
<ID>OUT</ID>162 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>260</ID>
<type>AE_SMALL_INVERTER</type>
<position>71.5,-31.5</position>
<input>
<ID>IN_0</ID>180 </input>
<output>
<ID>OUT_0</ID>181 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>227</ID>
<type>DA_FROM</type>
<position>149,-21.5</position>
<input>
<ID>IN_0</ID>22 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>228</ID>
<type>DA_FROM</type>
<position>150,-45.5</position>
<input>
<ID>IN_0</ID>20 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>229</ID>
<type>DA_FROM</type>
<position>150.5,-59.5</position>
<input>
<ID>IN_0</ID>19 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>230</ID>
<type>DA_FROM</type>
<position>148.5,-78</position>
<input>
<ID>IN_0</ID>23 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q4</lparam></gate>
<gate>
<ID>232</ID>
<type>AE_SMALL_INVERTER</type>
<position>66.5,-7.5</position>
<input>
<ID>IN_0</ID>154 </input>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>234</ID>
<type>AA_AND2</type>
<position>-22.5,-4</position>
<input>
<ID>IN_0</ID>167 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>127 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>240</ID>
<type>AE_SMALL_INVERTER</type>
<position>-17.5,-5</position>
<input>
<ID>IN_0</ID>155 </input>
<output>
<ID>OUT_0</ID>167 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>266</ID>
<type>DE_TO</type>
<position>185.5,-19</position>
<input>
<ID>IN_0</ID>187 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>241</ID>
<type>DE_TO</type>
<position>68.5,-15.5</position>
<input>
<ID>IN_0</ID>173 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>242</ID>
<type>DE_TO</type>
<position>68.5,-17.5</position>
<input>
<ID>IN_0</ID>169 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>243</ID>
<type>DE_TO</type>
<position>68.5,-19.5</position>
<input>
<ID>IN_0</ID>170 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>244</ID>
<type>DE_TO</type>
<position>67.5,-25</position>
<input>
<ID>IN_0</ID>179 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E</lparam></gate>
<gate>
<ID>245</ID>
<type>DE_TO</type>
<position>67.5,-27</position>
<input>
<ID>IN_0</ID>177 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>270</ID>
<type>DE_TO</type>
<position>185.5,-11</position>
<input>
<ID>IN_0</ID>183 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>246</ID>
<type>DE_TO</type>
<position>67.5,-29</position>
<input>
<ID>IN_0</ID>178 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>247</ID>
<type>DE_TO</type>
<position>68.5,-13.5</position>
<input>
<ID>IN_0</ID>168 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A</lparam></gate>
<gate>
<ID>264</ID>
<type>DE_TO</type>
<position>185.5,-15</position>
<input>
<ID>IN_0</ID>185 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C</lparam></gate>
<gate>
<ID>248</ID>
<type>DE_TO</type>
<position>67.5,-31.5</position>
<input>
<ID>IN_0</ID>180 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID H</lparam></gate>
<gate>
<ID>250</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-13.5</position>
<input>
<ID>IN_0</ID>168 </input>
<output>
<ID>OUT_0</ID>172 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>252</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-17.5</position>
<input>
<ID>IN_0</ID>169 </input>
<output>
<ID>OUT_0</ID>174 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>254</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-19.5</position>
<input>
<ID>IN_0</ID>170 </input>
<output>
<ID>OUT_0</ID>175 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>262</ID>
<type>EE_VDD</type>
<position>87,-11.5</position>
<output>
<ID>OUT_0</ID>182 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>265</ID>
<type>DE_TO</type>
<position>185.5,-17</position>
<input>
<ID>IN_0</ID>186 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D</lparam></gate>
<gate>
<ID>267</ID>
<type>DE_TO</type>
<position>185.5,-21</position>
<input>
<ID>IN_0</ID>188 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F</lparam></gate>
<gate>
<ID>268</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>201,-15.5</position>
<input>
<ID>IN_0</ID>183 </input>
<input>
<ID>IN_1</ID>184 </input>
<input>
<ID>IN_2</ID>185 </input>
<input>
<ID>IN_3</ID>186 </input>
<input>
<ID>IN_4</ID>187 </input>
<input>
<ID>IN_5</ID>188 </input>
<input>
<ID>IN_6</ID>189 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 114</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>269</ID>
<type>DE_TO</type>
<position>185.5,-23</position>
<input>
<ID>IN_0</ID>189 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>58,-38.5</position>
<input>
<ID>IN_0</ID>26 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>15</ID>
<type>AA_AND3</type>
<position>-21.5,-36.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>9 </input>
<input>
<ID>IN_2</ID>7 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>17</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16,-34.5</position>
<input>
<ID>IN_0</ID>29 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>18</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16,-36.5</position>
<input>
<ID>IN_0</ID>158 </input>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>67,-36</position>
<input>
<ID>IN_0</ID>157 </input>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>24</ID>
<type>DE_TO</type>
<position>-12.5,-38.5</position>
<input>
<ID>IN_0</ID>11 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>26</ID>
<type>DE_TO</type>
<position>68,-41</position>
<input>
<ID>IN_0</ID>57 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>27</ID>
<type>DE_TO</type>
<position>68,-43</position>
<input>
<ID>IN_0</ID>70 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>28</ID>
<type>DE_TO</type>
<position>68,-45</position>
<input>
<ID>IN_0</ID>69 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>30</ID>
<type>DE_TO</type>
<position>68,-50</position>
<input>
<ID>IN_0</ID>68 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E1</lparam></gate>
<gate>
<ID>32</ID>
<type>DE_TO</type>
<position>68,-52</position>
<input>
<ID>IN_0</ID>67 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F1</lparam></gate>
<gate>
<ID>37</ID>
<type>DE_TO</type>
<position>68,-54</position>
<input>
<ID>IN_0</ID>66 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G1</lparam></gate>
<gate>
<ID>39</ID>
<type>DE_TO</type>
<position>68.5,-38.5</position>
<input>
<ID>IN_0</ID>71 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>44</ID>
<type>DE_TO</type>
<position>68,-56.5</position>
<input>
<ID>IN_0</ID>65 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID H1</lparam></gate>
<gate>
<ID>46</ID>
<type>DE_TO</type>
<position>61,-47.5</position>
<input>
<ID>IN_0</ID>26 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>47</ID>
<type>DE_TO</type>
<position>80.5,-46</position>
<input>
<ID>IN_0</ID>27 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q1</lparam></gate>
<gate>
<ID>49</ID>
<type>DE_TO</type>
<position>185,-43</position>
<input>
<ID>IN_0</ID>46 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E1</lparam></gate>
<gate>
<ID>50</ID>
<type>DE_TO</type>
<position>185,-35</position>
<input>
<ID>IN_0</ID>34 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A1</lparam></gate>
<gate>
<ID>51</ID>
<type>DE_TO</type>
<position>185,-39</position>
<input>
<ID>IN_0</ID>37 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C1</lparam></gate>
<gate>
<ID>53</ID>
<type>DE_TO</type>
<position>185,-37</position>
<input>
<ID>IN_0</ID>36 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B1</lparam></gate>
<gate>
<ID>55</ID>
<type>DE_TO</type>
<position>185,-41</position>
<input>
<ID>IN_0</ID>44 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D1</lparam></gate>
<gate>
<ID>60</ID>
<type>DE_TO</type>
<position>185,-45</position>
<input>
<ID>IN_0</ID>47 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F1</lparam></gate>
<gate>
<ID>66</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>200.5,-39.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>36 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>44 </input>
<input>
<ID>IN_4</ID>46 </input>
<input>
<ID>IN_5</ID>47 </input>
<input>
<ID>IN_6</ID>54 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 2</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>67</ID>
<type>DE_TO</type>
<position>185,-47</position>
<input>
<ID>IN_0</ID>54 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G1</lparam></gate>
<gate>
<ID>69</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-37.5</position>
<input>
<ID>IN_0</ID>71 </input>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>76</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-41.5</position>
<input>
<ID>IN_0</ID>70 </input>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-43.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>85</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-50</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-52</position>
<input>
<ID>IN_0</ID>67 </input>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>89</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-54</position>
<input>
<ID>IN_0</ID>66 </input>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>91</ID>
<type>AE_SMALL_INVERTER</type>
<position>73.5,-56</position>
<input>
<ID>IN_0</ID>65 </input>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>93</ID>
<type>AA_AND3</type>
<position>-22,-66.5</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<input>
<ID>IN_2</ID>73 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>94</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16.5,-64.5</position>
<input>
<ID>IN_0</ID>160 </input>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>95</ID>
<type>AE_SMALL_INVERTER</type>
<position>-16.5,-66.5</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>74 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>96</ID>
<type>DE_TO</type>
<position>-13,-68.5</position>
<input>
<ID>IN_0</ID>75 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_AND2</type>
<position>53.5,-67.5</position>
<input>
<ID>IN_0</ID>83 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>98</ID>
<type>AE_SMALL_INVERTER</type>
<position>58.5,-66.5</position>
<input>
<ID>IN_0</ID>159 </input>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>99</ID>
<type>AA_AND3</type>
<position>-20,-97.5</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>78 </input>
<input>
<ID>IN_2</ID>77 </input>
<output>
<ID>OUT</ID>148 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>100</ID>
<type>AE_SMALL_INVERTER</type>
<position>-14.5,-95.5</position>
<input>
<ID>IN_0</ID>162 </input>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>101</ID>
<type>AE_SMALL_INVERTER</type>
<position>-14.5,-97.5</position>
<input>
<ID>IN_0</ID>49 </input>
<output>
<ID>OUT_0</ID>78 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>102</ID>
<type>DE_TO</type>
<position>-11,-99.5</position>
<input>
<ID>IN_0</ID>79 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_AND2</type>
<position>55.5,-98.5</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>80 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 180</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>104</ID>
<type>AE_SMALL_INVERTER</type>
<position>60.5,-97.5</position>
<input>
<ID>IN_0</ID>161 </input>
<output>
<ID>OUT_0</ID>80 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>105</ID>
<type>DE_TO</type>
<position>81.5,-71</position>
<input>
<ID>IN_0</ID>81 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>106</ID>
<type>DE_TO</type>
<position>85.5,-94</position>
<input>
<ID>IN_0</ID>82 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>107</ID>
<type>DE_TO</type>
<position>58.5,-68.5</position>
<input>
<ID>IN_0</ID>83 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q2</lparam></gate>
<gate>
<ID>108</ID>
<type>DE_TO</type>
<position>60.5,-99.5</position>
<input>
<ID>IN_0</ID>84 </input>
<gparam>angle 0.0</gparam>
<lparam>JUNCTION_ID Q3</lparam></gate>
<gate>
<ID>109</ID>
<type>DE_TO</type>
<position>68,-65.5</position>
<input>
<ID>IN_0</ID>98 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>110</ID>
<type>DE_TO</type>
<position>68,-67.5</position>
<input>
<ID>IN_0</ID>87 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>111</ID>
<type>DE_TO</type>
<position>68,-69.5</position>
<input>
<ID>IN_0</ID>88 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>112</ID>
<type>DE_TO</type>
<position>67.5,-74.5</position>
<input>
<ID>IN_0</ID>89 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E2</lparam></gate>
<gate>
<ID>113</ID>
<type>DE_TO</type>
<position>67.5,-76.5</position>
<input>
<ID>IN_0</ID>94 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F2</lparam></gate>
<gate>
<ID>114</ID>
<type>DE_TO</type>
<position>67.5,-78.5</position>
<input>
<ID>IN_0</ID>90 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G2</lparam></gate>
<gate>
<ID>115</ID>
<type>DE_TO</type>
<position>68.5,-63</position>
<input>
<ID>IN_0</ID>86 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>116</ID>
<type>DE_TO</type>
<position>67.5,-81</position>
<input>
<ID>IN_0</ID>91 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID H2</lparam></gate>
<gate>
<ID>117</ID>
<type>DE_TO</type>
<position>68,-87.5</position>
<input>
<ID>IN_0</ID>104 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>118</ID>
<type>DE_TO</type>
<position>68,-89.5</position>
<input>
<ID>IN_0</ID>171 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>119</ID>
<type>DE_TO</type>
<position>68,-91.5</position>
<input>
<ID>IN_0</ID>190 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>120</ID>
<type>DE_TO</type>
<position>68.5,-99</position>
<input>
<ID>IN_0</ID>103 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E3</lparam></gate>
<gate>
<ID>121</ID>
<type>DE_TO</type>
<position>68.5,-101</position>
<input>
<ID>IN_0</ID>106 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F3</lparam></gate>
<gate>
<ID>122</ID>
<type>DE_TO</type>
<position>68.5,-103</position>
<input>
<ID>IN_0</ID>193 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G3</lparam></gate>
<gate>
<ID>123</ID>
<type>DE_TO</type>
<position>68.5,-85</position>
<input>
<ID>IN_0</ID>101 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>124</ID>
<type>DE_TO</type>
<position>68.5,-105.5</position>
<input>
<ID>IN_0</ID>191 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID H3</lparam></gate>
<gate>
<ID>126</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-62</position>
<input>
<ID>IN_0</ID>86 </input>
<output>
<ID>OUT_0</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>128</ID>
<type>AE_SMALL_INVERTER</type>
<position>72,-67.5</position>
<input>
<ID>IN_0</ID>87 </input>
<output>
<ID>OUT_0</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>130</ID>
<type>AE_SMALL_INVERTER</type>
<position>72,-69.5</position>
<input>
<ID>IN_0</ID>88 </input>
<output>
<ID>OUT_0</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AE_SMALL_INVERTER</type>
<position>71.5,-74.5</position>
<input>
<ID>IN_0</ID>89 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>134</ID>
<type>AE_SMALL_INVERTER</type>
<position>71.5,-78.5</position>
<input>
<ID>IN_0</ID>90 </input>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>71.5,-81</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>146</ID>
<type>AE_SMALL_INVERTER</type>
<position>72,-87.5</position>
<input>
<ID>IN_0</ID>104 </input>
<output>
<ID>OUT_0</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>148</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-101</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>150</ID>
<type>DE_TO</type>
<position>183,-65.5</position>
<input>
<ID>IN_0</ID>123 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E2</lparam></gate>
<gate>
<ID>151</ID>
<type>DE_TO</type>
<position>183,-57.5</position>
<input>
<ID>IN_0</ID>119 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A2</lparam></gate>
<gate>
<ID>152</ID>
<type>DE_TO</type>
<position>183,-61.5</position>
<input>
<ID>IN_0</ID>121 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C2</lparam></gate>
<gate>
<ID>153</ID>
<type>DE_TO</type>
<position>183,-59.5</position>
<input>
<ID>IN_0</ID>120 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B2</lparam></gate>
<gate>
<ID>154</ID>
<type>DE_TO</type>
<position>183,-63.5</position>
<input>
<ID>IN_0</ID>122 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D2</lparam></gate>
<gate>
<ID>155</ID>
<type>DE_TO</type>
<position>183,-67.5</position>
<input>
<ID>IN_0</ID>124 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F2</lparam></gate>
<gate>
<ID>156</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>198.5,-62</position>
<input>
<ID>IN_0</ID>119 </input>
<input>
<ID>IN_1</ID>120 </input>
<input>
<ID>IN_2</ID>121 </input>
<input>
<ID>IN_3</ID>122 </input>
<input>
<ID>IN_4</ID>123 </input>
<input>
<ID>IN_5</ID>124 </input>
<input>
<ID>IN_6</ID>125 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 34</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>157</ID>
<type>DE_TO</type>
<position>183,-69.5</position>
<input>
<ID>IN_0</ID>125 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G2</lparam></gate>
<gate>
<ID>158</ID>
<type>DE_TO</type>
<position>182.5,-89.5</position>
<input>
<ID>IN_0</ID>116 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID E3</lparam></gate>
<gate>
<ID>159</ID>
<type>DE_TO</type>
<position>182.5,-81.5</position>
<input>
<ID>IN_0</ID>112 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID A3</lparam></gate>
<gate>
<ID>161</ID>
<type>DE_TO</type>
<position>182.5,-85.5</position>
<input>
<ID>IN_0</ID>114 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID C3</lparam></gate>
<gate>
<ID>162</ID>
<type>DE_TO</type>
<position>182.5,-83.5</position>
<input>
<ID>IN_0</ID>113 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B3</lparam></gate>
<gate>
<ID>163</ID>
<type>DE_TO</type>
<position>182.5,-87.5</position>
<input>
<ID>IN_0</ID>115 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID D3</lparam></gate>
<gate>
<ID>164</ID>
<type>DE_TO</type>
<position>182.5,-91.5</position>
<input>
<ID>IN_0</ID>117 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID F3</lparam></gate>
<gate>
<ID>205</ID>
<type>GI_LED_DISPLAY_8BIT</type>
<position>198,-86</position>
<input>
<ID>IN_0</ID>112 </input>
<input>
<ID>IN_1</ID>113 </input>
<input>
<ID>IN_2</ID>114 </input>
<input>
<ID>IN_3</ID>115 </input>
<input>
<ID>IN_4</ID>116 </input>
<input>
<ID>IN_5</ID>117 </input>
<input>
<ID>IN_6</ID>118 </input>
<gparam>VALUE_BOX -3.9,-3.9,3.9,4.9</gparam>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 89</lparam>
<lparam>INPUT_BITS 8</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_LOAD false</lparam>
<lparam>UNKNOWN_OUTPUTS false</lparam></gate>
<gate>
<ID>206</ID>
<type>DE_TO</type>
<position>182.5,-93.5</position>
<input>
<ID>IN_0</ID>118 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID G3</lparam></gate>
<gate>
<ID>207</ID>
<type>AE_SMALL_INVERTER</type>
<position>72,-89.5</position>
<input>
<ID>IN_0</ID>171 </input>
<output>
<ID>OUT_0</ID>176 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>208</ID>
<type>AE_SMALL_INVERTER</type>
<position>72.5,-105.5</position>
<input>
<ID>IN_0</ID>191 </input>
<output>
<ID>OUT_0</ID>192 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>210</ID>
<type>AA_LABEL</type>
<position>194,-3.5</position>
<gparam>LABEL_TEXT Nivel 1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>AA_LABEL</type>
<position>194,-29.5</position>
<gparam>LABEL_TEXT Nivel 2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>213</ID>
<type>AA_LABEL</type>
<position>194.5,-51.5</position>
<gparam>LABEL_TEXT Nivel 3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>215</ID>
<type>AA_LABEL</type>
<position>194,-74.5</position>
<gparam>LABEL_TEXT Nivel 4</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>-86,-17</position>
<gparam>LABEL_TEXT Contador 1</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>-87.5,-48.5</position>
<gparam>LABEL_TEXT Contador 2</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>-86.5,-75.5</position>
<gparam>LABEL_TEXT Contador 3</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_LABEL</type>
<position>-87,-107</position>
<gparam>LABEL_TEXT Contador 4</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>82</ID>
<type>EE_VDD</type>
<position>161.5,-46.5</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>263</ID>
<type>DE_TO</type>
<position>185.5,-13</position>
<input>
<ID>IN_0</ID>184 </input>
<gparam>angle 180</gparam>
<lparam>JUNCTION_ID B</lparam></gate>
<gate>
<ID>7</ID>
<type>AE_SMALL_INVERTER</type>
<position>-17.5,-3</position>
<input>
<ID>IN_0</ID>2 </input>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>angle 180</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>46.5,27</position>
<gparam>LABEL_TEXT Existem 2 conjuntos de 4 flip-flops em cada n�vel. O conjunto da direita eh o primeiro digito do numero e o da esquerda eh o segundo digito</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-19,15</position>
<gparam>LABEL_TEXT Quando o primeiro digito do nivel eh descoberto, o segundo comeca a ser contado</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-10,8</position>
<gparam>LABEL_TEXT Caso os dois digitos sejam descobertos, o nivel eh desbloqueado, partindo para o proximo</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>28,20.5</position>
<gparam>LABEL_TEXT Para a contagem comecar, o nivel anterior precisa estar desbloqueado. No caso do primeiro, ele comeca automaticamente</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>49 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-112,54,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-4,-103.5,54,-103.5</points>
<intersection>-4 149</intersection>
<intersection>1 23</intersection>
<intersection>12 21</intersection>
<intersection>22 19</intersection>
<intersection>33 12</intersection>
<intersection>43.5 5</intersection>
<intersection>52.5 151</intersection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>1,-112,55,-112</points>
<connection>
<GID>70</GID>
<name>J</name></connection>
<intersection>1 23</intersection>
<intersection>10.5 113</intersection>
<intersection>12 21</intersection>
<intersection>12.5 51</intersection>
<intersection>21 114</intersection>
<intersection>22 19</intersection>
<intersection>23.5 50</intersection>
<intersection>31.5 115</intersection>
<intersection>33 12</intersection>
<intersection>34 49</intersection>
<intersection>42 116</intersection>
<intersection>43.5 5</intersection>
<intersection>44.5 48</intersection>
<intersection>54 0</intersection>
<intersection>55 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-112,43.5,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>1,-108,55,-108</points>
<connection>
<GID>70</GID>
<name>K</name></connection>
<intersection>1 23</intersection>
<intersection>10.5 113</intersection>
<intersection>12 21</intersection>
<intersection>12.5 51</intersection>
<intersection>21 114</intersection>
<intersection>22 19</intersection>
<intersection>23.5 50</intersection>
<intersection>31.5 115</intersection>
<intersection>33 12</intersection>
<intersection>34 49</intersection>
<intersection>42 116</intersection>
<intersection>43.5 5</intersection>
<intersection>44.5 48</intersection>
<intersection>54 0</intersection>
<intersection>55 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>33,-112,33,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>22,-112,22,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>12,-112,12,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>1,-112,1,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>55,-112,55,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>44.5,-112,44.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>34,-112,34,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>23.5,-112,23.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>12.5,-112,12.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>10.5,-112,10.5,-108</points>
<connection>
<GID>74</GID>
<name>K</name></connection>
<connection>
<GID>74</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>21,-112,21,-108</points>
<connection>
<GID>73</GID>
<name>K</name></connection>
<connection>
<GID>73</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>31.5,-112,31.5,-108</points>
<connection>
<GID>72</GID>
<name>K</name></connection>
<connection>
<GID>72</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>42,-112,42,-108</points>
<connection>
<GID>71</GID>
<name>K</name></connection>
<connection>
<GID>71</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>149</ID>
<points>-4,-103.5,-4,-97.5</points>
<intersection>-103.5 1</intersection>
<intersection>-97.5 150</intersection></vsegment>
<hsegment>
<ID>150</ID>
<points>-12.5,-97.5,-4,-97.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-4 149</intersection></hsegment>
<vsegment>
<ID>151</ID>
<points>52.5,-103.5,52.5,-98.5</points>
<connection>
<GID>103</GID>
<name>OUT</name></connection>
<intersection>-103.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>51 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-112,23.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-110,23.5,-110</points>
<connection>
<GID>73</GID>
<name>clock</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-112,25.5,-112</points>
<connection>
<GID>72</GID>
<name>Q</name></connection>
<intersection>23.5 0</intersection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-117,25.5,-112</points>
<connection>
<GID>79</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment></shape></wire>
<wire>
<ID>52 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-112,12.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-110,12.5,-110</points>
<connection>
<GID>74</GID>
<name>clock</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-112,15,-112</points>
<connection>
<GID>73</GID>
<name>Q</name></connection>
<intersection>12.5 0</intersection>
<intersection>15 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-117,15,-112</points>
<intersection>-117 7</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>14.5,-117,15,-117</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment></shape></wire>
<wire>
<ID>8 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>34,-19,34,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>32,-17,34,-17</points>
<connection>
<GID>4</GID>
<name>clock</name></connection>
<intersection>34 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>34,-19,36.5,-19</points>
<connection>
<GID>2</GID>
<name>Q</name></connection>
<intersection>34 0</intersection>
<intersection>36.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36.5,-24,36.5,-19</points>
<intersection>-24 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>36,-24,36.5,-24</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>36.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>43 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>4,-86,4,-81</points>
<connection>
<GID>65</GID>
<name>IN_0</name></connection>
<connection>
<GID>59</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>2 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-19,54.5,-7.5</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection>
<intersection>-7.5 52</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2.5,-13,54.5,-13</points>
<intersection>2.5 23</intersection>
<intersection>12.5 21</intersection>
<intersection>22.5 19</intersection>
<intersection>33.5 12</intersection>
<intersection>44 5</intersection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2.5,-19,55.5,-19</points>
<connection>
<GID>1</GID>
<name>J</name></connection>
<connection>
<GID>2</GID>
<name>J</name></connection>
<connection>
<GID>4</GID>
<name>J</name></connection>
<connection>
<GID>5</GID>
<name>J</name></connection>
<connection>
<GID>6</GID>
<name>J</name></connection>
<intersection>2.5 23</intersection>
<intersection>12.5 21</intersection>
<intersection>13 51</intersection>
<intersection>22.5 19</intersection>
<intersection>24 50</intersection>
<intersection>33.5 12</intersection>
<intersection>34.5 49</intersection>
<intersection>44 5</intersection>
<intersection>45 48</intersection>
<intersection>54.5 0</intersection>
<intersection>55.5 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>44,-19,44,-12</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-13.5,-12,55.5,-12</points>
<intersection>-13.5 62</intersection>
<intersection>2.5 23</intersection>
<intersection>11 61</intersection>
<intersection>12.5 21</intersection>
<intersection>13 51</intersection>
<intersection>21.5 60</intersection>
<intersection>22.5 19</intersection>
<intersection>24 50</intersection>
<intersection>32 59</intersection>
<intersection>33.5 12</intersection>
<intersection>34.5 49</intersection>
<intersection>42.5 58</intersection>
<intersection>44 5</intersection>
<intersection>45 48</intersection>
<intersection>53 57</intersection>
<intersection>54.5 0</intersection>
<intersection>55.5 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>33.5,-19,33.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>22.5,-19,22.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>12.5,-19,12.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>2.5,-19,2.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-13 1</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>55.5,-19,55.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>45,-19,45,-12</points>
<intersection>-19 3</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>34.5,-19,34.5,-12</points>
<intersection>-19 3</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>24,-19,24,-12</points>
<intersection>-19 3</intersection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>13,-19,13,-12</points>
<intersection>-19 3</intersection>
<intersection>-12 7</intersection></vsegment>
<hsegment>
<ID>52</ID>
<points>54.5,-7.5,64.5,-7.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<vsegment>
<ID>57</ID>
<points>53,-15,53,-12</points>
<connection>
<GID>1</GID>
<name>K</name></connection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>58</ID>
<points>42.5,-15,42.5,-12</points>
<connection>
<GID>2</GID>
<name>K</name></connection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>59</ID>
<points>32,-15,32,-12</points>
<connection>
<GID>4</GID>
<name>K</name></connection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>60</ID>
<points>21.5,-15,21.5,-12</points>
<connection>
<GID>5</GID>
<name>K</name></connection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>61</ID>
<points>11,-15,11,-12</points>
<connection>
<GID>6</GID>
<name>K</name></connection>
<intersection>-12 7</intersection></vsegment>
<vsegment>
<ID>62</ID>
<points>-13.5,-12,-13.5,-3</points>
<intersection>-12 7</intersection>
<intersection>-3 63</intersection></vsegment>
<hsegment>
<ID>63</ID>
<points>-15.5,-3,-13.5,-3</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>-13.5 62</intersection></hsegment></shape></wire>
<wire>
<ID>1 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61.5,-23.5,61.5,-17</points>
<intersection>-23.5 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>53,-17,61.5,-17</points>
<connection>
<GID>1</GID>
<name>clock</name></connection>
<intersection>61.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-23.5,61.5,-23.5</points>
<connection>
<GID>3</GID>
<name>CLK</name></connection>
<intersection>61.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>3 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-19,46.5,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-17,46.5,-17</points>
<connection>
<GID>2</GID>
<name>clock</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46.5,-19,47,-19</points>
<connection>
<GID>1</GID>
<name>Q</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>53 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>4.5,-117,4.5,-112</points>
<connection>
<GID>81</GID>
<name>IN_0</name></connection>
<connection>
<GID>74</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>4 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>24,-19,24,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21.5,-17,24,-17</points>
<connection>
<GID>5</GID>
<name>clock</name></connection>
<intersection>24 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-19,26,-19</points>
<connection>
<GID>4</GID>
<name>Q</name></connection>
<intersection>24 0</intersection>
<intersection>26 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>26,-24,26,-19</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>-19 2</intersection></vsegment></shape></wire>
<wire>
<ID>5 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>13,-19,13,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>11,-17,13,-17</points>
<connection>
<GID>6</GID>
<name>clock</name></connection>
<intersection>13 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>13,-19,15.5,-19</points>
<connection>
<GID>5</GID>
<name>Q</name></connection>
<intersection>13 0</intersection>
<intersection>15.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15.5,-24,15.5,-19</points>
<intersection>-24 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>15,-24,15.5,-24</points>
<connection>
<GID>11</GID>
<name>IN_0</name></connection>
<intersection>15.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>48 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-116.5,61,-110</points>
<intersection>-116.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-110,61,-110</points>
<connection>
<GID>70</GID>
<name>clock</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58.5,-116.5,61,-116.5</points>
<connection>
<GID>77</GID>
<name>CLK</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>50 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-112,46,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-110,46,-110</points>
<connection>
<GID>71</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-112,46.5,-112</points>
<connection>
<GID>70</GID>
<name>Q</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>6 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>5,-24,5,-19</points>
<connection>
<GID>6</GID>
<name>Q</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147.5,-88.5,151.5,-88.5</points>
<intersection>147.5 5</intersection>
<intersection>151.5 6</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>147.5,-88.5,147.5,-80</points>
<intersection>-88.5 1</intersection>
<intersection>-80 7</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>151.5,-88.5,151.5,-80</points>
<intersection>-88.5 1</intersection>
<intersection>-80 8</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>144.5,-80,147.5,-80</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>146.5 10</intersection>
<intersection>147.5 5</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>151.5,-80,174.5,-80</points>
<connection>
<GID>13</GID>
<name>N_in0</name></connection>
<intersection>151.5 6</intersection></hsegment>
<vsegment>
<ID>10</ID>
<points>146.5,-80,146.5,-78</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>-80 7</intersection></vsegment></shape></wire>
<wire>
<ID>29 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-52,54,-38.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection>
<intersection>-38.5 133</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-43.5,54,-43.5</points>
<intersection>2 23</intersection>
<intersection>12 21</intersection>
<intersection>22 19</intersection>
<intersection>33 12</intersection>
<intersection>43.5 5</intersection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>2,-52,55,-52</points>
<connection>
<GID>19</GID>
<name>J</name></connection>
<intersection>2 23</intersection>
<intersection>10.5 113</intersection>
<intersection>12 21</intersection>
<intersection>12.5 51</intersection>
<intersection>21 114</intersection>
<intersection>22 19</intersection>
<intersection>23.5 50</intersection>
<intersection>31.5 115</intersection>
<intersection>33 12</intersection>
<intersection>34 49</intersection>
<intersection>42 116</intersection>
<intersection>43.5 5</intersection>
<intersection>44.5 48</intersection>
<intersection>54 0</intersection>
<intersection>55 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43.5,-52,43.5,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>2,-48,55,-48</points>
<connection>
<GID>19</GID>
<name>K</name></connection>
<intersection>2 23</intersection>
<intersection>10.5 113</intersection>
<intersection>12 21</intersection>
<intersection>12.5 51</intersection>
<intersection>21 114</intersection>
<intersection>22 19</intersection>
<intersection>23.5 50</intersection>
<intersection>31.5 115</intersection>
<intersection>33 12</intersection>
<intersection>34 49</intersection>
<intersection>42 116</intersection>
<intersection>43.5 5</intersection>
<intersection>44.5 48</intersection>
<intersection>54 0</intersection>
<intersection>55 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>33,-52,33,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>22,-52,22,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>12,-52,12,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>2,-52,2,-34.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection>
<intersection>-34.5 135</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>55,-52,55,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>44.5,-52,44.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>34,-52,34,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>23.5,-52,23.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>12.5,-52,12.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>10.5,-52,10.5,-48</points>
<connection>
<GID>25</GID>
<name>K</name></connection>
<connection>
<GID>25</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>21,-52,21,-48</points>
<connection>
<GID>52</GID>
<name>K</name></connection>
<connection>
<GID>52</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>31.5,-52,31.5,-48</points>
<connection>
<GID>23</GID>
<name>K</name></connection>
<connection>
<GID>23</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>42,-52,42,-48</points>
<connection>
<GID>21</GID>
<name>K</name></connection>
<connection>
<GID>21</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<hsegment>
<ID>133</ID>
<points>54,-38.5,55,-38.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>135</ID>
<points>-14,-34.5,2,-34.5</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>2 23</intersection></hsegment></shape></wire>
<wire>
<ID>28 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-56.5,61,-50</points>
<intersection>-56.5 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52.5,-50,61,-50</points>
<connection>
<GID>19</GID>
<name>clock</name></connection>
<intersection>61 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>57,-56.5,61,-56.5</points>
<connection>
<GID>29</GID>
<name>CLK</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>30 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46,-52,46,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-50,46,-50</points>
<connection>
<GID>21</GID>
<name>clock</name></connection>
<intersection>46 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>46,-52,46.5,-52</points>
<connection>
<GID>19</GID>
<name>Q</name></connection>
<intersection>46 0</intersection></hsegment></shape></wire>
<wire>
<ID>35 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-52,33.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-50,33.5,-50</points>
<connection>
<GID>23</GID>
<name>clock</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-52,36,-52</points>
<connection>
<GID>21</GID>
<name>Q</name></connection>
<intersection>33.5 0</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-57,36,-52</points>
<intersection>-57 5</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>35.5,-57,36,-57</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>31 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23.5,-52,23.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>21,-50,23.5,-50</points>
<connection>
<GID>52</GID>
<name>clock</name></connection>
<intersection>23.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23.5,-52,25.5,-52</points>
<connection>
<GID>23</GID>
<name>Q</name></connection>
<intersection>23.5 0</intersection>
<intersection>25.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25.5,-57,25.5,-52</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>-52 2</intersection></vsegment></shape></wire>
<wire>
<ID>32 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-52,12.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10.5,-50,12.5,-50</points>
<connection>
<GID>25</GID>
<name>clock</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12.5,-52,15,-52</points>
<connection>
<GID>52</GID>
<name>Q</name></connection>
<intersection>12.5 0</intersection>
<intersection>15 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>15,-57,15,-52</points>
<intersection>-57 5</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>14.5,-57,15,-57</points>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>15 3</intersection></hsegment></shape></wire>
<wire>
<ID>33 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>4.5,-57,4.5,-52</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<connection>
<GID>25</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>164 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116.5,-69.5,116.5,-61.5</points>
<intersection>-69.5 2</intersection>
<intersection>-61.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116.5,-61.5,139,-61.5</points>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>116.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-69.5,116.5,-69.5</points>
<connection>
<GID>221</GID>
<name>OUT</name></connection>
<intersection>116.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-86,156.5,-27.5</points>
<intersection>-86 17</intersection>
<intersection>-67.5 10</intersection>
<intersection>-51.5 4</intersection>
<intersection>-27.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>142.5,-27.5,156.5,-27.5</points>
<connection>
<GID>36</GID>
<name>clear</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>142.5,-51.5,161.5,-51.5</points>
<intersection>142.5 18</intersection>
<intersection>156.5 0</intersection>
<intersection>161.5 19</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>142,-67.5,156.5,-67.5</points>
<connection>
<GID>34</GID>
<name>clear</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>17</ID>
<points>141.5,-86,156.5,-86</points>
<connection>
<GID>45</GID>
<name>clear</name></connection>
<intersection>156.5 0</intersection></hsegment>
<vsegment>
<ID>18</ID>
<points>142.5,-51.5,142.5,-51</points>
<connection>
<GID>38</GID>
<name>clear</name></connection>
<intersection>-51.5 4</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>161.5,-51.5,161.5,-47.5</points>
<connection>
<GID>82</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>18 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>135,-32,139,-32</points>
<intersection>135 5</intersection>
<intersection>139 16</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>135,-83,135,-30.5</points>
<intersection>-83 21</intersection>
<intersection>-64.5 14</intersection>
<intersection>-48 12</intersection>
<intersection>-32 2</intersection>
<intersection>-30.5 27</intersection></vsegment>
<hsegment>
<ID>12</ID>
<points>135,-48,139.5,-48</points>
<connection>
<GID>38</GID>
<name>clock</name></connection>
<intersection>135 5</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>135,-64.5,139,-64.5</points>
<connection>
<GID>34</GID>
<name>clock</name></connection>
<intersection>135 5</intersection></hsegment>
<vsegment>
<ID>16</ID>
<points>139,-32,139,-24.5</points>
<intersection>-32 2</intersection>
<intersection>-24.5 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>139,-24.5,139.5,-24.5</points>
<connection>
<GID>36</GID>
<name>clock</name></connection>
<intersection>139 16</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>135,-83,138.5,-83</points>
<connection>
<GID>45</GID>
<name>clock</name></connection>
<intersection>135 5</intersection></hsegment>
<hsegment>
<ID>27</ID>
<points>132,-30.5,135,-30.5</points>
<connection>
<GID>160</GID>
<name>CLK</name></connection>
<intersection>135 5</intersection></hsegment></shape></wire>
<wire>
<ID>19 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>148,-71.5,151.5,-71.5</points>
<intersection>148 19</intersection>
<intersection>151.5 20</intersection></hsegment>
<vsegment>
<ID>19</ID>
<points>148,-71.5,148,-59.5</points>
<intersection>-71.5 2</intersection>
<intersection>-61.5 21</intersection>
<intersection>-59.5 24</intersection></vsegment>
<vsegment>
<ID>20</ID>
<points>151.5,-71.5,151.5,-61</points>
<intersection>-71.5 2</intersection>
<intersection>-61 22</intersection></vsegment>
<hsegment>
<ID>21</ID>
<points>145,-61.5,148,-61.5</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>148 19</intersection></hsegment>
<hsegment>
<ID>22</ID>
<points>151.5,-61,173.5,-61</points>
<connection>
<GID>40</GID>
<name>N_in0</name></connection>
<intersection>151.5 20</intersection></hsegment>
<hsegment>
<ID>24</ID>
<points>148,-59.5,148.5,-59.5</points>
<connection>
<GID>229</GID>
<name>IN_0</name></connection>
<intersection>148 19</intersection></hsegment></shape></wire>
<wire>
<ID>156 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>117,-21.5,117,-21</points>
<intersection>-21.5 1</intersection>
<intersection>-21 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>117,-21.5,139.5,-21.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>117 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94.5,-21,117,-21</points>
<connection>
<GID>214</GID>
<name>OUT</name></connection>
<intersection>117 0</intersection></hsegment></shape></wire>
<wire>
<ID>22 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>145.5,-15.5,151,-15.5</points>
<intersection>145.5 5</intersection>
<intersection>151 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>151,-17.5,151,-15.5</points>
<intersection>-17.5 8</intersection>
<intersection>-15.5 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>145.5,-21.5,145.5,-15.5</points>
<connection>
<GID>36</GID>
<name>OUT_0</name></connection>
<intersection>-21.5 12</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>151,-17.5,172,-17.5</points>
<connection>
<GID>41</GID>
<name>N_in0</name></connection>
<intersection>151 4</intersection></hsegment>
<hsegment>
<ID>12</ID>
<points>145.5,-21.5,147,-21.5</points>
<connection>
<GID>227</GID>
<name>IN_0</name></connection>
<intersection>145.5 5</intersection></hsegment></shape></wire>
<wire>
<ID>127 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-11.5,-19,-11.5,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-63.5,-13,-11.5,-13</points>
<intersection>-63.5 23</intersection>
<intersection>-53.5 21</intersection>
<intersection>-43.5 19</intersection>
<intersection>-32.5 12</intersection>
<intersection>-27 68</intersection>
<intersection>-22 5</intersection>
<intersection>-11.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-63.5,-19,-10.5,-19</points>
<connection>
<GID>165</GID>
<name>J</name></connection>
<connection>
<GID>166</GID>
<name>J</name></connection>
<connection>
<GID>168</GID>
<name>J</name></connection>
<connection>
<GID>169</GID>
<name>J</name></connection>
<connection>
<GID>170</GID>
<name>J</name></connection>
<intersection>-63.5 23</intersection>
<intersection>-53.5 21</intersection>
<intersection>-53 51</intersection>
<intersection>-43.5 19</intersection>
<intersection>-42 50</intersection>
<intersection>-32.5 12</intersection>
<intersection>-31.5 49</intersection>
<intersection>-22 5</intersection>
<intersection>-21 48</intersection>
<intersection>-11.5 0</intersection>
<intersection>-10.5 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-22,-19,-22,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-63.5,-15,-10.5,-15</points>
<connection>
<GID>165</GID>
<name>K</name></connection>
<connection>
<GID>166</GID>
<name>K</name></connection>
<connection>
<GID>168</GID>
<name>K</name></connection>
<connection>
<GID>169</GID>
<name>K</name></connection>
<connection>
<GID>170</GID>
<name>K</name></connection>
<intersection>-63.5 23</intersection>
<intersection>-53.5 21</intersection>
<intersection>-53 51</intersection>
<intersection>-43.5 19</intersection>
<intersection>-42 50</intersection>
<intersection>-32.5 12</intersection>
<intersection>-31.5 49</intersection>
<intersection>-22 5</intersection>
<intersection>-21 48</intersection>
<intersection>-11.5 0</intersection>
<intersection>-10.5 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-32.5,-19,-32.5,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-43.5,-19,-43.5,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-53.5,-19,-53.5,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-63.5,-19,-63.5,-13</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection>
<intersection>-13 1</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>-10.5,-19,-10.5,-15</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>-21,-19,-21,-15</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>-31.5,-19,-31.5,-15</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>-42,-19,-42,-15</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-53,-19,-53,-15</points>
<intersection>-19 3</intersection>
<intersection>-15 7</intersection></vsegment>
<vsegment>
<ID>68</ID>
<points>-27,-13,-27,-4</points>
<intersection>-13 1</intersection>
<intersection>-4 69</intersection></vsegment>
<hsegment>
<ID>69</ID>
<points>-27,-4,-25.5,-4</points>
<connection>
<GID>234</GID>
<name>OUT</name></connection>
<intersection>-27 68</intersection></hsegment></shape></wire>
<wire>
<ID>128 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-19,-19.5,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-23.5,-17,-19.5,-17</points>
<connection>
<GID>166</GID>
<name>clock</name></connection>
<intersection>-19.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-19.5,-19,-19,-19</points>
<connection>
<GID>165</GID>
<name>Q</name></connection>
<intersection>-19.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32,-19,-32,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34,-17,-32,-17</points>
<connection>
<GID>168</GID>
<name>clock</name></connection>
<intersection>-32 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32,-19,-29.5,-19</points>
<connection>
<GID>166</GID>
<name>Q</name></connection>
<intersection>-32 0</intersection>
<intersection>-29.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-29.5,-24,-29.5,-19</points>
<intersection>-24 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-30,-24,-29.5,-24</points>
<connection>
<GID>171</GID>
<name>IN_0</name></connection>
<intersection>-29.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>163 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>94.5,-45,139.5,-45</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<connection>
<GID>218</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>20 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>147,-54,156,-54</points>
<intersection>147 16</intersection>
<intersection>156 15</intersection></hsegment>
<vsegment>
<ID>15</ID>
<points>156,-54,156,-37.5</points>
<intersection>-54 1</intersection>
<intersection>-37.5 19</intersection></vsegment>
<vsegment>
<ID>16</ID>
<points>147,-54,147,-45</points>
<intersection>-54 1</intersection>
<intersection>-45.5 21</intersection>
<intersection>-45 18</intersection></vsegment>
<hsegment>
<ID>18</ID>
<points>145.5,-45,147,-45</points>
<connection>
<GID>38</GID>
<name>OUT_0</name></connection>
<intersection>147 16</intersection></hsegment>
<hsegment>
<ID>19</ID>
<points>156,-37.5,171,-37.5</points>
<connection>
<GID>43</GID>
<name>N_in0</name></connection>
<intersection>156 15</intersection></hsegment>
<hsegment>
<ID>21</ID>
<points>147,-45.5,148,-45.5</points>
<connection>
<GID>228</GID>
<name>IN_0</name></connection>
<intersection>147 16</intersection></hsegment></shape></wire>
<wire>
<ID>129 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42,-19,-42,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-44.5,-17,-42,-17</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<intersection>-42 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42,-19,-40,-19</points>
<connection>
<GID>168</GID>
<name>Q</name></connection>
<intersection>-42 0</intersection>
<intersection>-40 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40,-24,-40,-19</points>
<connection>
<GID>172</GID>
<name>IN_0</name></connection>
<intersection>-19 2</intersection></vsegment></shape></wire>
<wire>
<ID>130 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53,-19,-53,-17</points>
<intersection>-19 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55,-17,-53,-17</points>
<connection>
<GID>170</GID>
<name>clock</name></connection>
<intersection>-53 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53,-19,-50.5,-19</points>
<connection>
<GID>169</GID>
<name>Q</name></connection>
<intersection>-53 0</intersection>
<intersection>-50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-50.5,-24,-50.5,-19</points>
<intersection>-24 4</intersection>
<intersection>-19 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-51,-24,-50.5,-24</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-50.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>131 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-61,-24,-61,-19</points>
<connection>
<GID>174</GID>
<name>IN_0</name></connection>
<connection>
<GID>170</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>39 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>53.5,-81,53.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>0.5,-72.5,53.5,-72.5</points>
<intersection>0.5 23</intersection>
<intersection>11.5 21</intersection>
<intersection>21.5 19</intersection>
<intersection>32.5 12</intersection>
<intersection>43 5</intersection>
<intersection>50.5 133</intersection>
<intersection>53.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>0.5,-81,54.5,-81</points>
<connection>
<GID>42</GID>
<name>J</name></connection>
<intersection>0.5 23</intersection>
<intersection>10 113</intersection>
<intersection>11.5 21</intersection>
<intersection>12 51</intersection>
<intersection>20.5 114</intersection>
<intersection>21.5 19</intersection>
<intersection>23 50</intersection>
<intersection>31 115</intersection>
<intersection>32.5 12</intersection>
<intersection>33.5 49</intersection>
<intersection>41.5 116</intersection>
<intersection>43 5</intersection>
<intersection>44 48</intersection>
<intersection>53.5 0</intersection>
<intersection>54.5 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>43,-81,43,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>0.5,-77,54.5,-77</points>
<connection>
<GID>42</GID>
<name>K</name></connection>
<intersection>0.5 23</intersection>
<intersection>10 113</intersection>
<intersection>11.5 21</intersection>
<intersection>12 51</intersection>
<intersection>20.5 114</intersection>
<intersection>21.5 19</intersection>
<intersection>23 50</intersection>
<intersection>31 115</intersection>
<intersection>32.5 12</intersection>
<intersection>33.5 49</intersection>
<intersection>41.5 116</intersection>
<intersection>43 5</intersection>
<intersection>44 48</intersection>
<intersection>53.5 0</intersection>
<intersection>54.5 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>32.5,-81,32.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>21.5,-81,21.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>11.5,-81,11.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>0.5,-81,0.5,-66.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection>
<intersection>-66.5 135</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>54.5,-81,54.5,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>44,-81,44,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>33.5,-81,33.5,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>23,-81,23,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>12,-81,12,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>10,-81,10,-77</points>
<connection>
<GID>59</GID>
<name>K</name></connection>
<connection>
<GID>59</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>20.5,-81,20.5,-77</points>
<connection>
<GID>58</GID>
<name>K</name></connection>
<connection>
<GID>58</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>31,-81,31,-77</points>
<connection>
<GID>57</GID>
<name>K</name></connection>
<connection>
<GID>57</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>41.5,-81,41.5,-77</points>
<connection>
<GID>56</GID>
<name>K</name></connection>
<connection>
<GID>56</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>133</ID>
<points>50.5,-72.5,50.5,-67.5</points>
<connection>
<GID>97</GID>
<name>OUT</name></connection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>135</ID>
<points>-14.5,-66.5,0.5,-66.5</points>
<connection>
<GID>95</GID>
<name>IN_0</name></connection>
<intersection>0.5 23</intersection></hsegment></shape></wire>
<wire>
<ID>38 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-85.5,60.5,-79</points>
<intersection>-85.5 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>52,-79,60.5,-79</points>
<connection>
<GID>42</GID>
<name>clock</name></connection>
<intersection>60.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>58,-85.5,60.5,-85.5</points>
<connection>
<GID>61</GID>
<name>CLK</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45.5,-81,45.5,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-79,45.5,-79</points>
<connection>
<GID>56</GID>
<name>clock</name></connection>
<intersection>45.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>45.5,-81,46,-81</points>
<connection>
<GID>42</GID>
<name>Q</name></connection>
<intersection>45.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>165 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>116,-94,116,-80</points>
<intersection>-94 2</intersection>
<intersection>-80 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>116,-80,138.5,-80</points>
<connection>
<GID>45</GID>
<name>IN_0</name></connection>
<intersection>116 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-94,116,-94</points>
<connection>
<GID>224</GID>
<name>OUT</name></connection>
<intersection>116 0</intersection></hsegment></shape></wire>
<wire>
<ID>45 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-81,33,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-79,33,-79</points>
<connection>
<GID>57</GID>
<name>clock</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-81,35.5,-81</points>
<connection>
<GID>56</GID>
<name>Q</name></connection>
<intersection>33 0</intersection>
<intersection>35.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>35.5,-86,35.5,-81</points>
<intersection>-86 6</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>35,-86,35.5,-86</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>35.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>41 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-81,23,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-79,23,-79</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>23,-81,25,-81</points>
<connection>
<GID>57</GID>
<name>Q</name></connection>
<intersection>23 0</intersection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-86,25,-81</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>-81 2</intersection></vsegment></shape></wire>
<wire>
<ID>42 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12,-81,12,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>10,-79,12,-79</points>
<connection>
<GID>59</GID>
<name>clock</name></connection>
<intersection>12 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>12,-81,14.5,-81</points>
<connection>
<GID>58</GID>
<name>Q</name></connection>
<intersection>12 0</intersection>
<intersection>14.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>14.5,-86,14.5,-81</points>
<intersection>-86 6</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>14,-86,14.5,-86</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>14.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>55 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-112,33.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-110,33.5,-110</points>
<connection>
<GID>72</GID>
<name>clock</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-112,36,-112</points>
<connection>
<GID>71</GID>
<name>Q</name></connection>
<intersection>33.5 0</intersection>
<intersection>36 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-117,36,-112</points>
<intersection>-117 7</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>35.5,-117,36,-117</points>
<connection>
<GID>78</GID>
<name>IN_0</name></connection>
<intersection>36 3</intersection></hsegment></shape></wire>
<wire>
<ID>126 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-4.5,-23.5,-4.5,-17</points>
<intersection>-23.5 2</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13,-17,-4.5,-17</points>
<connection>
<GID>165</GID>
<name>clock</name></connection>
<intersection>-4.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-23.5,-4.5,-23.5</points>
<connection>
<GID>167</GID>
<name>CLK</name></connection>
<intersection>-4.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-52,-12,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-64,-43.5,-12,-43.5</points>
<intersection>-64 23</intersection>
<intersection>-54 21</intersection>
<intersection>-44 19</intersection>
<intersection>-33 12</intersection>
<intersection>-24.5 133</intersection>
<intersection>-22.5 5</intersection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-64,-52,-11,-52</points>
<connection>
<GID>175</GID>
<name>J</name></connection>
<intersection>-64 23</intersection>
<intersection>-55.5 113</intersection>
<intersection>-54 21</intersection>
<intersection>-53.5 51</intersection>
<intersection>-45 114</intersection>
<intersection>-44 19</intersection>
<intersection>-42.5 50</intersection>
<intersection>-34.5 115</intersection>
<intersection>-33 12</intersection>
<intersection>-32 49</intersection>
<intersection>-24 116</intersection>
<intersection>-22.5 5</intersection>
<intersection>-21.5 48</intersection>
<intersection>-12 0</intersection>
<intersection>-11 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-22.5,-52,-22.5,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-64,-48,-11,-48</points>
<connection>
<GID>175</GID>
<name>K</name></connection>
<intersection>-64 23</intersection>
<intersection>-55.5 113</intersection>
<intersection>-54 21</intersection>
<intersection>-53.5 51</intersection>
<intersection>-45 114</intersection>
<intersection>-44 19</intersection>
<intersection>-42.5 50</intersection>
<intersection>-34.5 115</intersection>
<intersection>-33 12</intersection>
<intersection>-32 49</intersection>
<intersection>-24 116</intersection>
<intersection>-22.5 5</intersection>
<intersection>-21.5 48</intersection>
<intersection>-12 0</intersection>
<intersection>-11 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-33,-52,-33,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-44,-52,-44,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-54,-52,-54,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-64,-52,-64,-43.5</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection>
<intersection>-43.5 1</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>-11,-52,-11,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>-21.5,-52,-21.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>-32,-52,-32,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>-42.5,-52,-42.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-53.5,-52,-53.5,-48</points>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>-55.5,-52,-55.5,-48</points>
<connection>
<GID>178</GID>
<name>K</name></connection>
<connection>
<GID>178</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>-45,-52,-45,-48</points>
<connection>
<GID>184</GID>
<name>K</name></connection>
<connection>
<GID>184</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>-34.5,-52,-34.5,-48</points>
<connection>
<GID>177</GID>
<name>K</name></connection>
<connection>
<GID>177</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-24,-52,-24,-48</points>
<connection>
<GID>176</GID>
<name>K</name></connection>
<connection>
<GID>176</GID>
<name>J</name></connection>
<intersection>-52 3</intersection>
<intersection>-48 7</intersection></vsegment>
<vsegment>
<ID>133</ID>
<points>-24.5,-43.5,-24.5,-36.5</points>
<connection>
<GID>15</GID>
<name>OUT</name></connection>
<intersection>-43.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>133 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-56.5,-5,-50</points>
<intersection>-56.5 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-50,-5,-50</points>
<connection>
<GID>175</GID>
<name>clock</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-9,-56.5,-5,-56.5</points>
<connection>
<GID>179</GID>
<name>CLK</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-52,-20,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-50,-20,-50</points>
<connection>
<GID>176</GID>
<name>clock</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20,-52,-19.5,-52</points>
<connection>
<GID>175</GID>
<name>Q</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>139 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-52,-32.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-50,-32.5,-50</points>
<connection>
<GID>177</GID>
<name>clock</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-52,-30,-52</points>
<connection>
<GID>176</GID>
<name>Q</name></connection>
<intersection>-32.5 0</intersection>
<intersection>-30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30,-57,-30,-52</points>
<intersection>-57 5</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-30.5,-57,-30,-57</points>
<connection>
<GID>185</GID>
<name>IN_0</name></connection>
<intersection>-30 3</intersection></hsegment></shape></wire>
<wire>
<ID>136 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-52,-42.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-50,-42.5,-50</points>
<connection>
<GID>184</GID>
<name>clock</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42.5,-52,-40.5,-52</points>
<connection>
<GID>177</GID>
<name>Q</name></connection>
<intersection>-42.5 0</intersection>
<intersection>-40.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40.5,-57,-40.5,-52</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>-52 2</intersection></vsegment></shape></wire>
<wire>
<ID>137 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-52,-53.5,-50</points>
<intersection>-52 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-50,-53.5,-50</points>
<connection>
<GID>178</GID>
<name>clock</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-52,-51,-52</points>
<connection>
<GID>184</GID>
<name>Q</name></connection>
<intersection>-53.5 0</intersection>
<intersection>-51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-51,-57,-51,-52</points>
<intersection>-57 5</intersection>
<intersection>-52 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-51.5,-57,-51,-57</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-51 3</intersection></hsegment></shape></wire>
<wire>
<ID>138 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-61.5,-57,-61.5,-52</points>
<connection>
<GID>182</GID>
<name>IN_0</name></connection>
<connection>
<GID>178</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>141 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12.5,-81,-12.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65.5,-72.5,-12.5,-72.5</points>
<intersection>-65.5 23</intersection>
<intersection>-54.5 21</intersection>
<intersection>-44.5 19</intersection>
<intersection>-33.5 12</intersection>
<intersection>-25 133</intersection>
<intersection>-23 5</intersection>
<intersection>-12.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-65.5,-81,-11.5,-81</points>
<connection>
<GID>183</GID>
<name>J</name></connection>
<intersection>-65.5 23</intersection>
<intersection>-56 113</intersection>
<intersection>-54.5 21</intersection>
<intersection>-54 51</intersection>
<intersection>-45.5 114</intersection>
<intersection>-44.5 19</intersection>
<intersection>-43 50</intersection>
<intersection>-35 115</intersection>
<intersection>-33.5 12</intersection>
<intersection>-32.5 49</intersection>
<intersection>-24.5 116</intersection>
<intersection>-23 5</intersection>
<intersection>-22 48</intersection>
<intersection>-12.5 0</intersection>
<intersection>-11.5 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-23,-81,-23,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-65.5,-77,-11.5,-77</points>
<connection>
<GID>183</GID>
<name>K</name></connection>
<intersection>-65.5 23</intersection>
<intersection>-56 113</intersection>
<intersection>-54.5 21</intersection>
<intersection>-54 51</intersection>
<intersection>-45.5 114</intersection>
<intersection>-44.5 19</intersection>
<intersection>-43 50</intersection>
<intersection>-35 115</intersection>
<intersection>-33.5 12</intersection>
<intersection>-32.5 49</intersection>
<intersection>-24.5 116</intersection>
<intersection>-23 5</intersection>
<intersection>-22 48</intersection>
<intersection>-12.5 0</intersection>
<intersection>-11.5 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-33.5,-81,-33.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-44.5,-81,-44.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-54.5,-81,-54.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-65.5,-81,-65.5,-72.5</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection>
<intersection>-72.5 1</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>-11.5,-81,-11.5,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>-22,-81,-22,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>-32.5,-81,-32.5,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>-43,-81,-43,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-54,-81,-54,-77</points>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>-56,-81,-56,-77</points>
<connection>
<GID>189</GID>
<name>K</name></connection>
<connection>
<GID>189</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>-45.5,-81,-45.5,-77</points>
<connection>
<GID>188</GID>
<name>K</name></connection>
<connection>
<GID>188</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>-35,-81,-35,-77</points>
<connection>
<GID>187</GID>
<name>K</name></connection>
<connection>
<GID>187</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-24.5,-81,-24.5,-77</points>
<connection>
<GID>186</GID>
<name>K</name></connection>
<connection>
<GID>186</GID>
<name>J</name></connection>
<intersection>-81 3</intersection>
<intersection>-77 7</intersection></vsegment>
<vsegment>
<ID>133</ID>
<points>-25,-72.5,-25,-66.5</points>
<connection>
<GID>93</GID>
<name>OUT</name></connection>
<intersection>-72.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>140 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5.5,-85.5,-5.5,-79</points>
<intersection>-85.5 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-14,-79,-5.5,-79</points>
<connection>
<GID>183</GID>
<name>clock</name></connection>
<intersection>-5.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8,-85.5,-5.5,-85.5</points>
<connection>
<GID>190</GID>
<name>CLK</name></connection>
<intersection>-5.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>142 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20.5,-81,-20.5,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24.5,-79,-20.5,-79</points>
<connection>
<GID>186</GID>
<name>clock</name></connection>
<intersection>-20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20.5,-81,-20,-81</points>
<connection>
<GID>183</GID>
<name>Q</name></connection>
<intersection>-20.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>146 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-33,-81,-33,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-35,-79,-33,-79</points>
<connection>
<GID>187</GID>
<name>clock</name></connection>
<intersection>-33 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-33,-81,-30.5,-81</points>
<connection>
<GID>186</GID>
<name>Q</name></connection>
<intersection>-33 0</intersection>
<intersection>-30.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30.5,-86,-30.5,-81</points>
<intersection>-86 6</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-31,-86,-30.5,-86</points>
<connection>
<GID>191</GID>
<name>IN_0</name></connection>
<intersection>-30.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>143 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-43,-81,-43,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45.5,-79,-43,-79</points>
<connection>
<GID>188</GID>
<name>clock</name></connection>
<intersection>-43 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-43,-81,-41,-81</points>
<connection>
<GID>187</GID>
<name>Q</name></connection>
<intersection>-43 0</intersection>
<intersection>-41 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-41,-86,-41,-81</points>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-81 2</intersection></vsegment></shape></wire>
<wire>
<ID>144 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-54,-81,-54,-79</points>
<intersection>-81 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-56,-79,-54,-79</points>
<connection>
<GID>189</GID>
<name>clock</name></connection>
<intersection>-54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-54,-81,-51.5,-81</points>
<connection>
<GID>188</GID>
<name>Q</name></connection>
<intersection>-54 0</intersection>
<intersection>-51.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-51.5,-86,-51.5,-81</points>
<intersection>-86 6</intersection>
<intersection>-81 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-52,-86,-51.5,-86</points>
<connection>
<GID>193</GID>
<name>IN_0</name></connection>
<intersection>-51.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>145 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-62,-86,-62,-81</points>
<connection>
<GID>194</GID>
<name>IN_0</name></connection>
<connection>
<GID>189</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>148 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-12,-112,-12,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-65,-103.5,-12,-103.5</points>
<intersection>-65 23</intersection>
<intersection>-54 21</intersection>
<intersection>-44 19</intersection>
<intersection>-33 12</intersection>
<intersection>-23 150</intersection>
<intersection>-22.5 5</intersection>
<intersection>-12 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-65,-112,-11,-112</points>
<connection>
<GID>195</GID>
<name>J</name></connection>
<intersection>-65 23</intersection>
<intersection>-55.5 113</intersection>
<intersection>-54 21</intersection>
<intersection>-53.5 51</intersection>
<intersection>-45 114</intersection>
<intersection>-44 19</intersection>
<intersection>-42.5 50</intersection>
<intersection>-34.5 115</intersection>
<intersection>-33 12</intersection>
<intersection>-32 49</intersection>
<intersection>-24 116</intersection>
<intersection>-22.5 5</intersection>
<intersection>-21.5 48</intersection>
<intersection>-12 0</intersection>
<intersection>-11 47</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-22.5,-112,-22.5,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-65,-108,-11,-108</points>
<connection>
<GID>195</GID>
<name>K</name></connection>
<intersection>-65 23</intersection>
<intersection>-55.5 113</intersection>
<intersection>-54 21</intersection>
<intersection>-53.5 51</intersection>
<intersection>-45 114</intersection>
<intersection>-44 19</intersection>
<intersection>-42.5 50</intersection>
<intersection>-34.5 115</intersection>
<intersection>-33 12</intersection>
<intersection>-32 49</intersection>
<intersection>-24 116</intersection>
<intersection>-22.5 5</intersection>
<intersection>-21.5 48</intersection>
<intersection>-12 0</intersection>
<intersection>-11 47</intersection></hsegment>
<vsegment>
<ID>12</ID>
<points>-33,-112,-33,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>19</ID>
<points>-44,-112,-44,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>21</ID>
<points>-54,-112,-54,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>23</ID>
<points>-65,-112,-65,-103.5</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection>
<intersection>-103.5 1</intersection></vsegment>
<vsegment>
<ID>47</ID>
<points>-11,-112,-11,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>48</ID>
<points>-21.5,-112,-21.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>49</ID>
<points>-32,-112,-32,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>50</ID>
<points>-42.5,-112,-42.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>51</ID>
<points>-53.5,-112,-53.5,-108</points>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>113</ID>
<points>-55.5,-112,-55.5,-108</points>
<connection>
<GID>199</GID>
<name>K</name></connection>
<connection>
<GID>199</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>114</ID>
<points>-45,-112,-45,-108</points>
<connection>
<GID>198</GID>
<name>K</name></connection>
<connection>
<GID>198</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>115</ID>
<points>-34.5,-112,-34.5,-108</points>
<connection>
<GID>197</GID>
<name>K</name></connection>
<connection>
<GID>197</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>116</ID>
<points>-24,-112,-24,-108</points>
<connection>
<GID>196</GID>
<name>K</name></connection>
<connection>
<GID>196</GID>
<name>J</name></connection>
<intersection>-112 3</intersection>
<intersection>-108 7</intersection></vsegment>
<vsegment>
<ID>150</ID>
<points>-23,-103.5,-23,-97.5</points>
<connection>
<GID>99</GID>
<name>OUT</name></connection>
<intersection>-103.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>147 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-5,-116.5,-5,-110</points>
<intersection>-116.5 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-13.5,-110,-5,-110</points>
<connection>
<GID>195</GID>
<name>clock</name></connection>
<intersection>-5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7.5,-116.5,-5,-116.5</points>
<connection>
<GID>200</GID>
<name>CLK</name></connection>
<intersection>-5 0</intersection></hsegment></shape></wire>
<wire>
<ID>149 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-20,-112,-20,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-24,-110,-20,-110</points>
<connection>
<GID>196</GID>
<name>clock</name></connection>
<intersection>-20 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-20,-112,-19.5,-112</points>
<connection>
<GID>195</GID>
<name>Q</name></connection>
<intersection>-20 0</intersection></hsegment></shape></wire>
<wire>
<ID>153 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-32.5,-112,-32.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-34.5,-110,-32.5,-110</points>
<connection>
<GID>197</GID>
<name>clock</name></connection>
<intersection>-32.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-32.5,-112,-30,-112</points>
<connection>
<GID>196</GID>
<name>Q</name></connection>
<intersection>-32.5 0</intersection>
<intersection>-30 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-30,-117,-30,-112</points>
<intersection>-117 7</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-30.5,-117,-30,-117</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-30 3</intersection></hsegment></shape></wire>
<wire>
<ID>150 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-42.5,-112,-42.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-45,-110,-42.5,-110</points>
<connection>
<GID>198</GID>
<name>clock</name></connection>
<intersection>-42.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-42.5,-112,-40.5,-112</points>
<connection>
<GID>197</GID>
<name>Q</name></connection>
<intersection>-42.5 0</intersection>
<intersection>-40.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-40.5,-117,-40.5,-112</points>
<connection>
<GID>202</GID>
<name>IN_0</name></connection>
<intersection>-112 2</intersection></vsegment></shape></wire>
<wire>
<ID>151 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-53.5,-112,-53.5,-110</points>
<intersection>-112 2</intersection>
<intersection>-110 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-55.5,-110,-53.5,-110</points>
<connection>
<GID>199</GID>
<name>clock</name></connection>
<intersection>-53.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-53.5,-112,-51,-112</points>
<connection>
<GID>198</GID>
<name>Q</name></connection>
<intersection>-53.5 0</intersection>
<intersection>-51 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-51,-117,-51,-112</points>
<intersection>-117 7</intersection>
<intersection>-112 2</intersection></vsegment>
<hsegment>
<ID>7</ID>
<points>-51.5,-117,-51,-117</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-51 3</intersection></hsegment></shape></wire>
<wire>
<ID>152 </ID>
<shape>
<vsegment>
<ID>3</ID>
<points>-61.5,-117,-61.5,-112</points>
<connection>
<GID>204</GID>
<name>IN_0</name></connection>
<connection>
<GID>199</GID>
<name>Q</name></connection></vsegment></shape></wire>
<wire>
<ID>172 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-13.5,76,-13.5</points>
<connection>
<GID>212</GID>
<name>IN_0</name></connection>
<connection>
<GID>250</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>173 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-15.5,76,-15.5</points>
<connection>
<GID>212</GID>
<name>IN_1</name></connection>
<connection>
<GID>241</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>174 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-17.5,76,-17.5</points>
<connection>
<GID>212</GID>
<name>IN_2</name></connection>
<connection>
<GID>252</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>175 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-19.5,76,-19.5</points>
<connection>
<GID>212</GID>
<name>IN_3</name></connection>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>154 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-19,85,-16.5</points>
<intersection>-19 1</intersection>
<intersection>-16.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-19,88.5,-19</points>
<connection>
<GID>214</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82,-16.5,85,-16.5</points>
<connection>
<GID>212</GID>
<name>OUT</name></connection>
<intersection>82.5 3</intersection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>82.5,-16.5,82.5,-7.5</points>
<intersection>-16.5 2</intersection>
<intersection>-7.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>68.5,-7.5,82.5,-7.5</points>
<connection>
<GID>232</GID>
<name>IN_0</name></connection>
<intersection>82.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>182 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>87,-21,87,-12.5</points>
<connection>
<GID>262</GID>
<name>OUT_0</name></connection>
<intersection>-21 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>87,-21,88.5,-21</points>
<connection>
<GID>214</GID>
<name>IN_1</name></connection>
<intersection>87 0</intersection></hsegment></shape></wire>
<wire>
<ID>155 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-29,85,-23</points>
<intersection>-29 2</intersection>
<intersection>-23 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-23,88.5,-23</points>
<connection>
<GID>214</GID>
<name>IN_2</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-29,85,-29</points>
<connection>
<GID>216</GID>
<name>OUT</name></connection>
<intersection>84 3</intersection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>84,-29,84,-5</points>
<intersection>-29 2</intersection>
<intersection>-5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-15.5,-5,84,-5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>84 3</intersection></hsegment></shape></wire>
<wire>
<ID>179 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-26,73,-25</points>
<intersection>-26 1</intersection>
<intersection>-25 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-26,75.5,-26</points>
<connection>
<GID>216</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-25,73,-25</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>177 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-28,73,-27</points>
<intersection>-28 1</intersection>
<intersection>-27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-28,75.5,-28</points>
<connection>
<GID>216</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-27,73,-27</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>178 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-30,73,-29</points>
<intersection>-30 1</intersection>
<intersection>-29 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-30,75.5,-30</points>
<connection>
<GID>216</GID>
<name>IN_2</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69.5,-29,73,-29</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>181 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-32,75,-31.5</points>
<intersection>-32 1</intersection>
<intersection>-31.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-32,75.5,-32</points>
<connection>
<GID>216</GID>
<name>IN_3</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-31.5,75,-31.5</points>
<connection>
<GID>260</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>58 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-37.5,76,-37.5</points>
<connection>
<GID>217</GID>
<name>IN_0</name></connection>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>57 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-41,73,-39.5</points>
<intersection>-41 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-39.5,76,-39.5</points>
<connection>
<GID>217</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-41,73,-41</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>59 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-41.5,76,-41.5</points>
<connection>
<GID>217</GID>
<name>IN_2</name></connection>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>60 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75.5,-43.5,76,-43.5</points>
<connection>
<GID>217</GID>
<name>IN_3</name></connection>
<connection>
<GID>83</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>157 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-43,85,-36</points>
<intersection>-43 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-43,88.5,-43</points>
<connection>
<GID>218</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>69,-36,85,-36</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<intersection>82 4</intersection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>82,-40.5,82,-36</points>
<connection>
<GID>217</GID>
<name>OUT</name></connection>
<intersection>-36 2</intersection></vsegment></shape></wire>
<wire>
<ID>27 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-46,88.5,-45</points>
<connection>
<GID>218</GID>
<name>IN_1</name></connection>
<intersection>-46 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>82.5,-46,88.5,-46</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>158 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-53,85,-47</points>
<intersection>-53 2</intersection>
<intersection>-47 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-47,88.5,-47</points>
<connection>
<GID>218</GID>
<name>IN_2</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81.5,-53,85,-53</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>83.5 3</intersection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>83.5,-53,83.5,-33.5</points>
<intersection>-53 2</intersection>
<intersection>-33.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-11,-33.5,83.5,-33.5</points>
<intersection>-11 5</intersection>
<intersection>83.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-11,-36.5,-11,-33.5</points>
<intersection>-36.5 6</intersection>
<intersection>-33.5 4</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-14,-36.5,-11,-36.5</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-11 5</intersection></hsegment></shape></wire>
<wire>
<ID>61 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-50,75.5,-50</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>62 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-52,75.5,-52</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>63 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-54,75.5,-54</points>
<connection>
<GID>219</GID>
<name>IN_2</name></connection>
<connection>
<GID>89</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>64 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-56,75.5,-56</points>
<connection>
<GID>219</GID>
<name>IN_3</name></connection>
<connection>
<GID>91</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>99 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-62,76,-62</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>98 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-65.5,73,-64</points>
<intersection>-65.5 2</intersection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-64,76,-64</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-65.5,73,-65.5</points>
<connection>
<GID>109</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>97 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-67.5,75,-66</points>
<intersection>-67.5 2</intersection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-66,76,-66</points>
<connection>
<GID>220</GID>
<name>IN_2</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-67.5,75,-67.5</points>
<connection>
<GID>128</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>96 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-69.5,75,-68</points>
<intersection>-69.5 2</intersection>
<intersection>-68 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-68,76,-68</points>
<connection>
<GID>220</GID>
<name>IN_3</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-69.5,75,-69.5</points>
<connection>
<GID>130</GID>
<name>OUT_0</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>159 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-67.5,85,-58.5</points>
<intersection>-67.5 1</intersection>
<intersection>-65 6</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-67.5,88.5,-67.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>60.5,-58.5,85,-58.5</points>
<intersection>60.5 4</intersection>
<intersection>85 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>60.5,-66.5,60.5,-58.5</points>
<connection>
<GID>98</GID>
<name>IN_0</name></connection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>82,-65,85,-65</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>81 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88.5,-71,88.5,-69.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>-71 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>83.5,-71,88.5,-71</points>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>88.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>160 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-77.5,84.5,-60</points>
<intersection>-77.5 5</intersection>
<intersection>-71.5 1</intersection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-71.5,88.5,-71.5</points>
<connection>
<GID>221</GID>
<name>IN_2</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-14.5,-60,84.5,-60</points>
<intersection>-14.5 3</intersection>
<intersection>84.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-14.5,-64.5,-14.5,-60</points>
<connection>
<GID>94</GID>
<name>IN_0</name></connection>
<intersection>-60 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>81.5,-77.5,84.5,-77.5</points>
<connection>
<GID>222</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-74.5,75.5,-74.5</points>
<connection>
<GID>222</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>94 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-76.5,75.5,-76.5</points>
<connection>
<GID>222</GID>
<name>IN_1</name></connection>
<connection>
<GID>113</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>93 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>73.5,-78.5,75.5,-78.5</points>
<connection>
<GID>222</GID>
<name>IN_2</name></connection>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>92 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-81,74.5,-80.5</points>
<intersection>-81 2</intersection>
<intersection>-80.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-80.5,75.5,-80.5</points>
<connection>
<GID>222</GID>
<name>IN_3</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-81,74.5,-81</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>101 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>73,-86.5,73,-85</points>
<intersection>-86.5 1</intersection>
<intersection>-85 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>73,-86.5,75.5,-86.5</points>
<connection>
<GID>223</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70.5,-85,73,-85</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>73 0</intersection></hsegment></shape></wire>
<wire>
<ID>108 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-88.5,74.5,-87.5</points>
<intersection>-88.5 1</intersection>
<intersection>-87.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-88.5,75.5,-88.5</points>
<connection>
<GID>223</GID>
<name>IN_1</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-87.5,74.5,-87.5</points>
<connection>
<GID>146</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>176 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-90.5,74.5,-89.5</points>
<intersection>-90.5 1</intersection>
<intersection>-89.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-90.5,75.5,-90.5</points>
<connection>
<GID>223</GID>
<name>IN_2</name></connection>
<intersection>74.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-89.5,74.5,-89.5</points>
<connection>
<GID>207</GID>
<name>OUT_0</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>190 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>72.5,-92.5,72.5,-91.5</points>
<intersection>-92.5 1</intersection>
<intersection>-91.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>72.5,-92.5,75.5,-92.5</points>
<connection>
<GID>223</GID>
<name>IN_3</name></connection>
<intersection>72.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-91.5,72.5,-91.5</points>
<connection>
<GID>119</GID>
<name>IN_0</name></connection>
<intersection>72.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>161 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-92,84.5,-83.5</points>
<intersection>-92 1</intersection>
<intersection>-89.5 5</intersection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-92,88,-92</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>62.5,-83.5,84.5,-83.5</points>
<intersection>62.5 3</intersection>
<intersection>84.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>62.5,-97.5,62.5,-83.5</points>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>81.5,-89.5,84.5,-89.5</points>
<connection>
<GID>223</GID>
<name>OUT</name></connection>
<intersection>84.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>82 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>87.5,-94,88,-94</points>
<connection>
<GID>224</GID>
<name>IN_1</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>162 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84.5,-107,84.5,-96</points>
<intersection>-107 2</intersection>
<intersection>-96 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84.5,-96,88,-96</points>
<connection>
<GID>224</GID>
<name>IN_2</name></connection>
<intersection>84.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-7,-107,84.5,-107</points>
<intersection>-7 5</intersection>
<intersection>81 4</intersection>
<intersection>84.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>81,-107,81,-102</points>
<connection>
<GID>225</GID>
<name>OUT</name></connection>
<intersection>-107 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-7,-107,-7,-95.5</points>
<intersection>-107 2</intersection>
<intersection>-95.5 6</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-12.5,-95.5,-7,-95.5</points>
<connection>
<GID>100</GID>
<name>IN_0</name></connection>
<intersection>-7 5</intersection></hsegment></shape></wire>
<wire>
<ID>103 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-99,75,-99</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<connection>
<GID>120</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>110 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>74.5,-101,75,-101</points>
<connection>
<GID>225</GID>
<name>IN_1</name></connection>
<connection>
<GID>148</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>193 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70.5,-103,75,-103</points>
<connection>
<GID>225</GID>
<name>IN_2</name></connection>
<connection>
<GID>122</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>192 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>74.5,-105.5,74.5,-105</points>
<connection>
<GID>208</GID>
<name>OUT_0</name></connection>
<intersection>-105 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>74.5,-105,75,-105</points>
<connection>
<GID>225</GID>
<name>IN_3</name></connection>
<intersection>74.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>180 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-31.5,69.5,-31.5</points>
<connection>
<GID>260</GID>
<name>IN_0</name></connection>
<connection>
<GID>248</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>167 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-5,-19.5,-5</points>
<connection>
<GID>234</GID>
<name>IN_0</name></connection>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>12 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-19.5,-3,-19.5,-3</points>
<connection>
<GID>234</GID>
<name>IN_1</name></connection>
<connection>
<GID>7</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>187 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-19,191.5,-14.5</points>
<intersection>-19 2</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-14.5,196,-14.5</points>
<connection>
<GID>268</GID>
<name>IN_4</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-19,191.5,-19</points>
<connection>
<GID>266</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>169 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-17.5,70.5,-17.5</points>
<connection>
<GID>242</GID>
<name>IN_0</name></connection>
<connection>
<GID>252</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>170 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-19.5,70.5,-19.5</points>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<connection>
<GID>254</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>183 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-18.5,191.5,-11</points>
<intersection>-18.5 6</intersection>
<intersection>-11 5</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>187.5,-11,191.5,-11</points>
<connection>
<GID>270</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>191.5,-18.5,196,-18.5</points>
<connection>
<GID>268</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>185 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-16.5,191.5,-15</points>
<intersection>-16.5 4</intersection>
<intersection>-15 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-15,191.5,-15</points>
<connection>
<GID>264</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>191.5,-16.5,196,-16.5</points>
<connection>
<GID>268</GID>
<name>IN_2</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>168 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-13.5,70.5,-13.5</points>
<connection>
<GID>247</GID>
<name>IN_0</name></connection>
<connection>
<GID>250</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>186 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-17,191.5,-15.5</points>
<intersection>-17 2</intersection>
<intersection>-15.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-15.5,196,-15.5</points>
<connection>
<GID>268</GID>
<name>IN_3</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-17,191.5,-17</points>
<connection>
<GID>265</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>188 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-21,191.5,-13.5</points>
<intersection>-21 2</intersection>
<intersection>-13.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-13.5,196,-13.5</points>
<connection>
<GID>268</GID>
<name>IN_5</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-21,191.5,-21</points>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>184 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-17.5,191.5,-13</points>
<intersection>-17.5 4</intersection>
<intersection>-13 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187.5,-13,191.5,-13</points>
<connection>
<GID>263</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>191.5,-17.5,196,-17.5</points>
<connection>
<GID>268</GID>
<name>IN_1</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>189 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191.5,-23,191.5,-12.5</points>
<intersection>-23 2</intersection>
<intersection>-12.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191.5,-12.5,196,-12.5</points>
<connection>
<GID>268</GID>
<name>IN_6</name></connection>
<intersection>191.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187.5,-23,191.5,-23</points>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>191.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-47.5,61,-39.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>59,-47.5,61,-47.5</points>
<connection>
<GID>46</GID>
<name>IN_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>10 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>61,-37.5,61,-36</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>-36 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>61,-36,65,-36</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>61 0</intersection></hsegment></shape></wire>
<wire>
<ID>11 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18.5,-38.5,-14.5,-38.5</points>
<connection>
<GID>15</GID>
<name>IN_0</name></connection>
<connection>
<GID>24</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18.5,-36.5,-18,-36.5</points>
<connection>
<GID>15</GID>
<name>IN_1</name></connection>
<connection>
<GID>18</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-18.5,-34.5,-18,-34.5</points>
<connection>
<GID>15</GID>
<name>IN_2</name></connection>
<connection>
<GID>17</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>70 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-43,70.5,-41.5</points>
<intersection>-43 2</intersection>
<intersection>-41.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-41.5,71.5,-41.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-43,70.5,-43</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>69 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-45,70.5,-43.5</points>
<intersection>-45 2</intersection>
<intersection>-43.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-43.5,71.5,-43.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-45,70.5,-45</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>68 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-50,71.5,-50</points>
<connection>
<GID>85</GID>
<name>IN_0</name></connection>
<connection>
<GID>30</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>67 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-52,71.5,-52</points>
<connection>
<GID>87</GID>
<name>IN_0</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>66 </ID>
<shape>
<hsegment>
<ID>2</ID>
<points>70,-54,71.5,-54</points>
<connection>
<GID>89</GID>
<name>IN_0</name></connection>
<connection>
<GID>37</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>71 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-38.5,70.5,-37.5</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70.5,-37.5,71.5,-37.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>70.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>71,-56.5,71,-56</points>
<intersection>-56.5 2</intersection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>71,-56,71.5,-56</points>
<connection>
<GID>91</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>70,-56.5,71,-56.5</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>71 0</intersection></hsegment></shape></wire>
<wire>
<ID>46 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-43,191,-38.5</points>
<intersection>-43 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-38.5,195.5,-38.5</points>
<connection>
<GID>66</GID>
<name>IN_4</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-43,191,-43</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>34 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-42.5,191,-35</points>
<intersection>-42.5 4</intersection>
<intersection>-35 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>187,-35,191,-35</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>191,-42.5,195.5,-42.5</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>37 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-40.5,191,-39</points>
<intersection>-40.5 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-40.5,195.5,-40.5</points>
<connection>
<GID>66</GID>
<name>IN_2</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-39,191,-39</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>36 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-41.5,191,-37</points>
<intersection>-41.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-41.5,195.5,-41.5</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-37,191,-37</points>
<connection>
<GID>53</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>44 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-41,191,-39.5</points>
<intersection>-41 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-39.5,195.5,-39.5</points>
<connection>
<GID>66</GID>
<name>IN_3</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-41,191,-41</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>47 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-45,191,-37.5</points>
<intersection>-45 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-37.5,195.5,-37.5</points>
<connection>
<GID>66</GID>
<name>IN_5</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-45,191,-45</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>54 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>191,-47,191,-36.5</points>
<intersection>-47 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>191,-36.5,195.5,-36.5</points>
<connection>
<GID>66</GID>
<name>IN_6</name></connection>
<intersection>191 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>187,-47,191,-47</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>191 0</intersection></hsegment></shape></wire>
<wire>
<ID>75 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-68.5,-15,-68.5</points>
<connection>
<GID>93</GID>
<name>IN_0</name></connection>
<connection>
<GID>96</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>74 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-66.5,-18.5,-66.5</points>
<connection>
<GID>95</GID>
<name>OUT_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>73 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-19,-64.5,-18.5,-64.5</points>
<connection>
<GID>94</GID>
<name>OUT_0</name></connection>
<connection>
<GID>93</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>83 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-68.5,56.5,-68.5</points>
<connection>
<GID>97</GID>
<name>IN_0</name></connection>
<connection>
<GID>107</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>76 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-66.5,56.5,-66.5</points>
<connection>
<GID>97</GID>
<name>IN_1</name></connection>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>79 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-99.5,-13,-99.5</points>
<connection>
<GID>99</GID>
<name>IN_0</name></connection>
<connection>
<GID>102</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>78 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-97.5,-16.5,-97.5</points>
<connection>
<GID>101</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>77 </ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-17,-95.5,-16.5,-95.5</points>
<connection>
<GID>100</GID>
<name>OUT_0</name></connection>
<connection>
<GID>99</GID>
<name>IN_2</name></connection></hsegment></shape></wire>
<wire>
<ID>84 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-99.5,58.5,-99.5</points>
<connection>
<GID>103</GID>
<name>IN_0</name></connection>
<connection>
<GID>108</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>80 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>58.5,-97.5,58.5,-97.5</points>
<connection>
<GID>103</GID>
<name>IN_1</name></connection>
<connection>
<GID>104</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>87 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-67.5,70,-67.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<connection>
<GID>128</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>88 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-69.5,70,-69.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<connection>
<GID>130</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>89 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-74.5,69.5,-74.5</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<connection>
<GID>132</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>90 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-78.5,69.5,-78.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<connection>
<GID>134</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>86 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-63,70.5,-62</points>
<connection>
<GID>126</GID>
<name>IN_0</name></connection>
<connection>
<GID>115</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>91 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-81,69.5,-81</points>
<connection>
<GID>116</GID>
<name>IN_0</name></connection>
<connection>
<GID>136</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>104 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-87.5,70,-87.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<connection>
<GID>146</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>171 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-89.5,70,-89.5</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<connection>
<GID>207</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>106 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-101,70.5,-101</points>
<connection>
<GID>121</GID>
<name>IN_0</name></connection>
<connection>
<GID>148</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>191 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70.5,-105.5,70.5,-105.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<connection>
<GID>208</GID>
<name>IN_0</name></connection></vsegment></shape></wire>
<wire>
<ID>123 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-65.5,189,-61</points>
<intersection>-65.5 2</intersection>
<intersection>-61 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-61,193.5,-61</points>
<connection>
<GID>156</GID>
<name>IN_4</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-65.5,189,-65.5</points>
<connection>
<GID>150</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>119 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-65,189,-57.5</points>
<intersection>-65 4</intersection>
<intersection>-57.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>185,-57.5,189,-57.5</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>189,-65,193.5,-65</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>121 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-63,189,-61.5</points>
<intersection>-63 1</intersection>
<intersection>-61.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-63,193.5,-63</points>
<connection>
<GID>156</GID>
<name>IN_2</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-61.5,189,-61.5</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>120 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-64,189,-59.5</points>
<intersection>-64 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-64,193.5,-64</points>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-59.5,189,-59.5</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>122 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-63.5,189,-62</points>
<intersection>-63.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-62,193.5,-62</points>
<connection>
<GID>156</GID>
<name>IN_3</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-63.5,189,-63.5</points>
<connection>
<GID>154</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>124 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-67.5,189,-60</points>
<intersection>-67.5 2</intersection>
<intersection>-60 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-60,193.5,-60</points>
<connection>
<GID>156</GID>
<name>IN_5</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-67.5,189,-67.5</points>
<connection>
<GID>155</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>125 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>189,-69.5,189,-59</points>
<intersection>-69.5 2</intersection>
<intersection>-59 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>189,-59,193.5,-59</points>
<connection>
<GID>156</GID>
<name>IN_6</name></connection>
<intersection>189 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>185,-69.5,189,-69.5</points>
<connection>
<GID>157</GID>
<name>IN_0</name></connection>
<intersection>189 0</intersection></hsegment></shape></wire>
<wire>
<ID>116 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-89.5,188.5,-85</points>
<intersection>-89.5 2</intersection>
<intersection>-85 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-85,193,-85</points>
<connection>
<GID>205</GID>
<name>IN_4</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-89.5,188.5,-89.5</points>
<connection>
<GID>158</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>112 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-89,188.5,-81.5</points>
<intersection>-89 4</intersection>
<intersection>-81.5 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>184.5,-81.5,188.5,-81.5</points>
<connection>
<GID>159</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>188.5,-89,193,-89</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>114 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-87,188.5,-85.5</points>
<intersection>-87 1</intersection>
<intersection>-85.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-87,193,-87</points>
<connection>
<GID>205</GID>
<name>IN_2</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-85.5,188.5,-85.5</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>113 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-88,188.5,-83.5</points>
<intersection>-88 1</intersection>
<intersection>-83.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-88,193,-88</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-83.5,188.5,-83.5</points>
<connection>
<GID>162</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>115 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-87.5,188.5,-86</points>
<intersection>-87.5 2</intersection>
<intersection>-86 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-86,193,-86</points>
<connection>
<GID>205</GID>
<name>IN_3</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-87.5,188.5,-87.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>117 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-91.5,188.5,-84</points>
<intersection>-91.5 2</intersection>
<intersection>-84 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-84,193,-84</points>
<connection>
<GID>205</GID>
<name>IN_5</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-91.5,188.5,-91.5</points>
<connection>
<GID>164</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>118 </ID>
<shape>
<vsegment>
<ID>0</ID>
<points>188.5,-93.5,188.5,-83</points>
<intersection>-93.5 2</intersection>
<intersection>-83 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>188.5,-83,193,-83</points>
<connection>
<GID>205</GID>
<name>IN_6</name></connection>
<intersection>188.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>184.5,-93.5,188.5,-93.5</points>
<connection>
<GID>206</GID>
<name>IN_0</name></connection>
<intersection>188.5 0</intersection></hsegment></shape></wire></page 0></circuit>